module dadda16(out_end,out, a, b);

	input [15:0]a;
	input [15:0]b;
	output [15:0]out;
	output out_end;
 

 /************************** AND gate DOT PRODUCT matrix ********************************/ 
	wire P_0_0;
	and A_0_0(P_0_0, a[0], b[0]);
	wire P_0_1;
	and A_0_1(P_0_1, a[0], b[1]);
	wire P_0_2;
	and A_0_2(P_0_2, a[0], b[2]);
	wire P_0_3;
	and A_0_3(P_0_3, a[0], b[3]);
	wire P_0_4;
	and A_0_4(P_0_4, a[0], b[4]);
	wire P_0_5;
	and A_0_5(P_0_5, a[0], b[5]);
	wire P_0_6;
	and A_0_6(P_0_6, a[0], b[6]);
	wire P_0_7;
	and A_0_7(P_0_7, a[0], b[7]);
	wire P_0_8;
	and A_0_8(P_0_8, a[0], b[8]);
	wire P_0_9;
	and A_0_9(P_0_9, a[0], b[9]);
	wire P_0_10;
	and A_0_10(P_0_10, a[0], b[10]);
	wire P_0_11;
	and A_0_11(P_0_11, a[0], b[11]);
	wire P_0_12;
	and A_0_12(P_0_12, a[0], b[12]);
	wire P_0_13;
	and A_0_13(P_0_13, a[0], b[13]);
	wire P_0_14;
	and A_0_14(P_0_14, a[0], b[14]);
	wire P_0_15;
	and A_0_15(P_0_15, a[0], b[15]);
	wire P_1_0;
	and A_1_0(P_1_0, a[1], b[0]);
	wire P_1_1;
	and A_1_1(P_1_1, a[1], b[1]);
	wire P_1_2;
	and A_1_2(P_1_2, a[1], b[2]);
	wire P_1_3;
	and A_1_3(P_1_3, a[1], b[3]);
	wire P_1_4;
	and A_1_4(P_1_4, a[1], b[4]);
	wire P_1_5;
	and A_1_5(P_1_5, a[1], b[5]);
	wire P_1_6;
	and A_1_6(P_1_6, a[1], b[6]);
	wire P_1_7;
	and A_1_7(P_1_7, a[1], b[7]);
	wire P_1_8;
	and A_1_8(P_1_8, a[1], b[8]);
	wire P_1_9;
	and A_1_9(P_1_9, a[1], b[9]);
	wire P_1_10;
	and A_1_10(P_1_10, a[1], b[10]);
	wire P_1_11;
	and A_1_11(P_1_11, a[1], b[11]);
	wire P_1_12;
	and A_1_12(P_1_12, a[1], b[12]);
	wire P_1_13;
	and A_1_13(P_1_13, a[1], b[13]);
	wire P_1_14;
	and A_1_14(P_1_14, a[1], b[14]);
	wire P_1_15;
	and A_1_15(P_1_15, a[1], b[15]);
	wire P_2_0;
	and A_2_0(P_2_0, a[2], b[0]);
	wire P_2_1;
	and A_2_1(P_2_1, a[2], b[1]);
	wire P_2_2;
	and A_2_2(P_2_2, a[2], b[2]);
	wire P_2_3;
	and A_2_3(P_2_3, a[2], b[3]);
	wire P_2_4;
	and A_2_4(P_2_4, a[2], b[4]);
	wire P_2_5;
	and A_2_5(P_2_5, a[2], b[5]);
	wire P_2_6;
	and A_2_6(P_2_6, a[2], b[6]);
	wire P_2_7;
	and A_2_7(P_2_7, a[2], b[7]);
	wire P_2_8;
	and A_2_8(P_2_8, a[2], b[8]);
	wire P_2_9;
	and A_2_9(P_2_9, a[2], b[9]);
	wire P_2_10;
	and A_2_10(P_2_10, a[2], b[10]);
	wire P_2_11;
	and A_2_11(P_2_11, a[2], b[11]);
	wire P_2_12;
	and A_2_12(P_2_12, a[2], b[12]);
	wire P_2_13;
	and A_2_13(P_2_13, a[2], b[13]);
	wire P_2_14;
	and A_2_14(P_2_14, a[2], b[14]);
	wire P_2_15;
	and A_2_15(P_2_15, a[2], b[15]);
	wire P_3_0;
	and A_3_0(P_3_0, a[3], b[0]);
	wire P_3_1;
	and A_3_1(P_3_1, a[3], b[1]);
	wire P_3_2;
	and A_3_2(P_3_2, a[3], b[2]);
	wire P_3_3;
	and A_3_3(P_3_3, a[3], b[3]);
	wire P_3_4;
	and A_3_4(P_3_4, a[3], b[4]);
	wire P_3_5;
	and A_3_5(P_3_5, a[3], b[5]);
	wire P_3_6;
	and A_3_6(P_3_6, a[3], b[6]);
	wire P_3_7;
	and A_3_7(P_3_7, a[3], b[7]);
	wire P_3_8;
	and A_3_8(P_3_8, a[3], b[8]);
	wire P_3_9;
	and A_3_9(P_3_9, a[3], b[9]);
	wire P_3_10;
	and A_3_10(P_3_10, a[3], b[10]);
	wire P_3_11;
	and A_3_11(P_3_11, a[3], b[11]);
	wire P_3_12;
	and A_3_12(P_3_12, a[3], b[12]);
	wire P_3_13;
	and A_3_13(P_3_13, a[3], b[13]);
	wire P_3_14;
	and A_3_14(P_3_14, a[3], b[14]);
	wire P_3_15;
	and A_3_15(P_3_15, a[3], b[15]);
	wire P_4_0;
	and A_4_0(P_4_0, a[4], b[0]);
	wire P_4_1;
	and A_4_1(P_4_1, a[4], b[1]);
	wire P_4_2;
	and A_4_2(P_4_2, a[4], b[2]);
	wire P_4_3;
	and A_4_3(P_4_3, a[4], b[3]);
	wire P_4_4;
	and A_4_4(P_4_4, a[4], b[4]);
	wire P_4_5;
	and A_4_5(P_4_5, a[4], b[5]);
	wire P_4_6;
	and A_4_6(P_4_6, a[4], b[6]);
	wire P_4_7;
	and A_4_7(P_4_7, a[4], b[7]);
	wire P_4_8;
	and A_4_8(P_4_8, a[4], b[8]);
	wire P_4_9;
	and A_4_9(P_4_9, a[4], b[9]);
	wire P_4_10;
	and A_4_10(P_4_10, a[4], b[10]);
	wire P_4_11;
	and A_4_11(P_4_11, a[4], b[11]);
	wire P_4_12;
	and A_4_12(P_4_12, a[4], b[12]);
	wire P_4_13;
	and A_4_13(P_4_13, a[4], b[13]);
	wire P_4_14;
	and A_4_14(P_4_14, a[4], b[14]);
	wire P_4_15;
	and A_4_15(P_4_15, a[4], b[15]);
	wire P_5_0;
	and A_5_0(P_5_0, a[5], b[0]);
	wire P_5_1;
	and A_5_1(P_5_1, a[5], b[1]);
	wire P_5_2;
	and A_5_2(P_5_2, a[5], b[2]);
	wire P_5_3;
	and A_5_3(P_5_3, a[5], b[3]);
	wire P_5_4;
	and A_5_4(P_5_4, a[5], b[4]);
	wire P_5_5;
	and A_5_5(P_5_5, a[5], b[5]);
	wire P_5_6;
	and A_5_6(P_5_6, a[5], b[6]);
	wire P_5_7;
	and A_5_7(P_5_7, a[5], b[7]);
	wire P_5_8;
	and A_5_8(P_5_8, a[5], b[8]);
	wire P_5_9;
	and A_5_9(P_5_9, a[5], b[9]);
	wire P_5_10;
	and A_5_10(P_5_10, a[5], b[10]);
	wire P_5_11;
	and A_5_11(P_5_11, a[5], b[11]);
	wire P_5_12;
	and A_5_12(P_5_12, a[5], b[12]);
	wire P_5_13;
	and A_5_13(P_5_13, a[5], b[13]);
	wire P_5_14;
	and A_5_14(P_5_14, a[5], b[14]);
	wire P_5_15;
	and A_5_15(P_5_15, a[5], b[15]);
	wire P_6_0;
	and A_6_0(P_6_0, a[6], b[0]);
	wire P_6_1;
	and A_6_1(P_6_1, a[6], b[1]);
	wire P_6_2;
	and A_6_2(P_6_2, a[6], b[2]);
	wire P_6_3;
	and A_6_3(P_6_3, a[6], b[3]);
	wire P_6_4;
	and A_6_4(P_6_4, a[6], b[4]);
	wire P_6_5;
	and A_6_5(P_6_5, a[6], b[5]);
	wire P_6_6;
	and A_6_6(P_6_6, a[6], b[6]);
	wire P_6_7;
	and A_6_7(P_6_7, a[6], b[7]);
	wire P_6_8;
	and A_6_8(P_6_8, a[6], b[8]);
	wire P_6_9;
	and A_6_9(P_6_9, a[6], b[9]);
	wire P_6_10;
	and A_6_10(P_6_10, a[6], b[10]);
	wire P_6_11;
	and A_6_11(P_6_11, a[6], b[11]);
	wire P_6_12;
	and A_6_12(P_6_12, a[6], b[12]);
	wire P_6_13;
	and A_6_13(P_6_13, a[6], b[13]);
	wire P_6_14;
	and A_6_14(P_6_14, a[6], b[14]);
	wire P_6_15;
	and A_6_15(P_6_15, a[6], b[15]);
	wire P_7_0;
	and A_7_0(P_7_0, a[7], b[0]);
	wire P_7_1;
	and A_7_1(P_7_1, a[7], b[1]);
	wire P_7_2;
	and A_7_2(P_7_2, a[7], b[2]);
	wire P_7_3;
	and A_7_3(P_7_3, a[7], b[3]);
	wire P_7_4;
	and A_7_4(P_7_4, a[7], b[4]);
	wire P_7_5;
	and A_7_5(P_7_5, a[7], b[5]);
	wire P_7_6;
	and A_7_6(P_7_6, a[7], b[6]);
	wire P_7_7;
	and A_7_7(P_7_7, a[7], b[7]);
	wire P_7_8;
	and A_7_8(P_7_8, a[7], b[8]);
	wire P_7_9;
	and A_7_9(P_7_9, a[7], b[9]);
	wire P_7_10;
	and A_7_10(P_7_10, a[7], b[10]);
	wire P_7_11;
	and A_7_11(P_7_11, a[7], b[11]);
	wire P_7_12;
	and A_7_12(P_7_12, a[7], b[12]);
	wire P_7_13;
	and A_7_13(P_7_13, a[7], b[13]);
	wire P_7_14;
	and A_7_14(P_7_14, a[7], b[14]);
	wire P_7_15;
	and A_7_15(P_7_15, a[7], b[15]);
	wire P_8_0;
	and A_8_0(P_8_0, a[8], b[0]);
	wire P_8_1;
	and A_8_1(P_8_1, a[8], b[1]);
	wire P_8_2;
	and A_8_2(P_8_2, a[8], b[2]);
	wire P_8_3;
	and A_8_3(P_8_3, a[8], b[3]);
	wire P_8_4;
	and A_8_4(P_8_4, a[8], b[4]);
	wire P_8_5;
	and A_8_5(P_8_5, a[8], b[5]);
	wire P_8_6;
	and A_8_6(P_8_6, a[8], b[6]);
	wire P_8_7;
	and A_8_7(P_8_7, a[8], b[7]);
	wire P_8_8;
	and A_8_8(P_8_8, a[8], b[8]);
	wire P_8_9;
	and A_8_9(P_8_9, a[8], b[9]);
	wire P_8_10;
	and A_8_10(P_8_10, a[8], b[10]);
	wire P_8_11;
	and A_8_11(P_8_11, a[8], b[11]);
	wire P_8_12;
	and A_8_12(P_8_12, a[8], b[12]);
	wire P_8_13;
	and A_8_13(P_8_13, a[8], b[13]);
	wire P_8_14;
	and A_8_14(P_8_14, a[8], b[14]);
	wire P_8_15;
	and A_8_15(P_8_15, a[8], b[15]);
	wire P_9_0;
	and A_9_0(P_9_0, a[9], b[0]);
	wire P_9_1;
	and A_9_1(P_9_1, a[9], b[1]);
	wire P_9_2;
	and A_9_2(P_9_2, a[9], b[2]);
	wire P_9_3;
	and A_9_3(P_9_3, a[9], b[3]);
	wire P_9_4;
	and A_9_4(P_9_4, a[9], b[4]);
	wire P_9_5;
	and A_9_5(P_9_5, a[9], b[5]);
	wire P_9_6;
	and A_9_6(P_9_6, a[9], b[6]);
	wire P_9_7;
	and A_9_7(P_9_7, a[9], b[7]);
	wire P_9_8;
	and A_9_8(P_9_8, a[9], b[8]);
	wire P_9_9;
	and A_9_9(P_9_9, a[9], b[9]);
	wire P_9_10;
	and A_9_10(P_9_10, a[9], b[10]);
	wire P_9_11;
	and A_9_11(P_9_11, a[9], b[11]);
	wire P_9_12;
	and A_9_12(P_9_12, a[9], b[12]);
	wire P_9_13;
	and A_9_13(P_9_13, a[9], b[13]);
	wire P_9_14;
	and A_9_14(P_9_14, a[9], b[14]);
	wire P_9_15;
	and A_9_15(P_9_15, a[9], b[15]);
	wire P_10_0;
	and A_10_0(P_10_0, a[10], b[0]);
	wire P_10_1;
	and A_10_1(P_10_1, a[10], b[1]);
	wire P_10_2;
	and A_10_2(P_10_2, a[10], b[2]);
	wire P_10_3;
	and A_10_3(P_10_3, a[10], b[3]);
	wire P_10_4;
	and A_10_4(P_10_4, a[10], b[4]);
	wire P_10_5;
	and A_10_5(P_10_5, a[10], b[5]);
	wire P_10_6;
	and A_10_6(P_10_6, a[10], b[6]);
	wire P_10_7;
	and A_10_7(P_10_7, a[10], b[7]);
	wire P_10_8;
	and A_10_8(P_10_8, a[10], b[8]);
	wire P_10_9;
	and A_10_9(P_10_9, a[10], b[9]);
	wire P_10_10;
	and A_10_10(P_10_10, a[10], b[10]);
	wire P_10_11;
	and A_10_11(P_10_11, a[10], b[11]);
	wire P_10_12;
	and A_10_12(P_10_12, a[10], b[12]);
	wire P_10_13;
	and A_10_13(P_10_13, a[10], b[13]);
	wire P_10_14;
	and A_10_14(P_10_14, a[10], b[14]);
	wire P_10_15;
	and A_10_15(P_10_15, a[10], b[15]);
	wire P_11_0;
	and A_11_0(P_11_0, a[11], b[0]);
	wire P_11_1;
	and A_11_1(P_11_1, a[11], b[1]);
	wire P_11_2;
	and A_11_2(P_11_2, a[11], b[2]);
	wire P_11_3;
	and A_11_3(P_11_3, a[11], b[3]);
	wire P_11_4;
	and A_11_4(P_11_4, a[11], b[4]);
	wire P_11_5;
	and A_11_5(P_11_5, a[11], b[5]);
	wire P_11_6;
	and A_11_6(P_11_6, a[11], b[6]);
	wire P_11_7;
	and A_11_7(P_11_7, a[11], b[7]);
	wire P_11_8;
	and A_11_8(P_11_8, a[11], b[8]);
	wire P_11_9;
	and A_11_9(P_11_9, a[11], b[9]);
	wire P_11_10;
	and A_11_10(P_11_10, a[11], b[10]);
	wire P_11_11;
	and A_11_11(P_11_11, a[11], b[11]);
	wire P_11_12;
	and A_11_12(P_11_12, a[11], b[12]);
	wire P_11_13;
	and A_11_13(P_11_13, a[11], b[13]);
	wire P_11_14;
	and A_11_14(P_11_14, a[11], b[14]);
	wire P_11_15;
	and A_11_15(P_11_15, a[11], b[15]);
	wire P_12_0;
	and A_12_0(P_12_0, a[12], b[0]);
	wire P_12_1;
	and A_12_1(P_12_1, a[12], b[1]);
	wire P_12_2;
	and A_12_2(P_12_2, a[12], b[2]);
	wire P_12_3;
	and A_12_3(P_12_3, a[12], b[3]);
	wire P_12_4;
	and A_12_4(P_12_4, a[12], b[4]);
	wire P_12_5;
	and A_12_5(P_12_5, a[12], b[5]);
	wire P_12_6;
	and A_12_6(P_12_6, a[12], b[6]);
	wire P_12_7;
	and A_12_7(P_12_7, a[12], b[7]);
	wire P_12_8;
	and A_12_8(P_12_8, a[12], b[8]);
	wire P_12_9;
	and A_12_9(P_12_9, a[12], b[9]);
	wire P_12_10;
	and A_12_10(P_12_10, a[12], b[10]);
	wire P_12_11;
	and A_12_11(P_12_11, a[12], b[11]);
	wire P_12_12;
	and A_12_12(P_12_12, a[12], b[12]);
	wire P_12_13;
	and A_12_13(P_12_13, a[12], b[13]);
	wire P_12_14;
	and A_12_14(P_12_14, a[12], b[14]);
	wire P_12_15;
	and A_12_15(P_12_15, a[12], b[15]);
	wire P_13_0;
	and A_13_0(P_13_0, a[13], b[0]);
	wire P_13_1;
	and A_13_1(P_13_1, a[13], b[1]);
	wire P_13_2;
	and A_13_2(P_13_2, a[13], b[2]);
	wire P_13_3;
	and A_13_3(P_13_3, a[13], b[3]);
	wire P_13_4;
	and A_13_4(P_13_4, a[13], b[4]);
	wire P_13_5;
	and A_13_5(P_13_5, a[13], b[5]);
	wire P_13_6;
	and A_13_6(P_13_6, a[13], b[6]);
	wire P_13_7;
	and A_13_7(P_13_7, a[13], b[7]);
	wire P_13_8;
	and A_13_8(P_13_8, a[13], b[8]);
	wire P_13_9;
	and A_13_9(P_13_9, a[13], b[9]);
	wire P_13_10;
	and A_13_10(P_13_10, a[13], b[10]);
	wire P_13_11;
	and A_13_11(P_13_11, a[13], b[11]);
	wire P_13_12;
	and A_13_12(P_13_12, a[13], b[12]);
	wire P_13_13;
	and A_13_13(P_13_13, a[13], b[13]);
	wire P_13_14;
	and A_13_14(P_13_14, a[13], b[14]);
	wire P_13_15;
	and A_13_15(P_13_15, a[13], b[15]);
	wire P_14_0;
	and A_14_0(P_14_0, a[14], b[0]);
	wire P_14_1;
	and A_14_1(P_14_1, a[14], b[1]);
	wire P_14_2;
	and A_14_2(P_14_2, a[14], b[2]);
	wire P_14_3;
	and A_14_3(P_14_3, a[14], b[3]);
	wire P_14_4;
	and A_14_4(P_14_4, a[14], b[4]);
	wire P_14_5;
	and A_14_5(P_14_5, a[14], b[5]);
	wire P_14_6;
	and A_14_6(P_14_6, a[14], b[6]);
	wire P_14_7;
	and A_14_7(P_14_7, a[14], b[7]);
	wire P_14_8;
	and A_14_8(P_14_8, a[14], b[8]);
	wire P_14_9;
	and A_14_9(P_14_9, a[14], b[9]);
	wire P_14_10;
	and A_14_10(P_14_10, a[14], b[10]);
	wire P_14_11;
	and A_14_11(P_14_11, a[14], b[11]);
	wire P_14_12;
	and A_14_12(P_14_12, a[14], b[12]);
	wire P_14_13;
	and A_14_13(P_14_13, a[14], b[13]);
	wire P_14_14;
	and A_14_14(P_14_14, a[14], b[14]);
	wire P_14_15;
	and A_14_15(P_14_15, a[14], b[15]);
	wire P_15_0;
	and A_15_0(P_15_0, a[15], b[0]);
	wire P_15_1;
	and A_15_1(P_15_1, a[15], b[1]);
	wire P_15_2;
	and A_15_2(P_15_2, a[15], b[2]);
	wire P_15_3;
	and A_15_3(P_15_3, a[15], b[3]);
	wire P_15_4;
	and A_15_4(P_15_4, a[15], b[4]);
	wire P_15_5;
	and A_15_5(P_15_5, a[15], b[5]);
	wire P_15_6;
	and A_15_6(P_15_6, a[15], b[6]);
	wire P_15_7;
	and A_15_7(P_15_7, a[15], b[7]);
	wire P_15_8;
	and A_15_8(P_15_8, a[15], b[8]);
	wire P_15_9;
	and A_15_9(P_15_9, a[15], b[9]);
	wire P_15_10;
	and A_15_10(P_15_10, a[15], b[10]);
	wire P_15_11;
	and A_15_11(P_15_11, a[15], b[11]);
	wire P_15_12;
	and A_15_12(P_15_12, a[15], b[12]);
	wire P_15_13;
	and A_15_13(P_15_13, a[15], b[13]);
	wire P_15_14;
	and A_15_14(P_15_14, a[15], b[14]);
	wire P_15_15;
	and A_15_15(P_15_15, a[15], b[15]);
 

	wire [2:0] cout1;
	wire [2:0] cout2;
	wire [2:0] cout3;
	wire [2:0] cout4;
	wire [2:0] cout5;
	wire [2:0] cout6;
	wire [2:0] cout7;
	wire [2:0] cout8;
	wire [2:0] cout9;
	wire [2:0] cout10;
	wire [2:0] cout11;
	wire [2:0] cout12;
	wire [2:0] cout13;
	wire [2:0] cout14;
	wire [2:0] cout15;
	wire [2:0] cout16;
	wire [2:0] cout17;
	wire [2:0] cout18;
	wire [2:0] cout19;
	wire [2:0] cout20;
	wire [2:0] cout21;

	wire gout1;
	wire gout2;
	wire gout3;
	wire gout4;
	wire gout5;
	wire gout6;
	wire gout7;
	wire gout8;
	wire gout9;
	wire gout10;
	wire gout11;
	wire gout12;
	wire gout13;
	wire gout14;
	wire gout15;
	wire gout16;
	wire gout17;
	wire gout18;
	wire gout19;
	wire gout20;
	wire gout21;

	wire pout1;
	wire pout2;
	wire pout3;
	wire pout4;
	wire pout5;
	wire pout6;
	wire pout7;
	wire pout8;
	wire pout9;
	wire pout10;
	wire pout11;
	wire pout12;
	wire pout13;
	wire pout14;
	wire pout15;
	wire pout16;
	wire pout17;
	wire pout18;
	wire pout19;
	wire pout20;
	wire pout21;

	wire [3:0] la1;
	wire [3:0] lb1;
	wire [3:0] la2;
	wire [3:0] lb2;
	wire [3:0] la3;
	wire [3:0] lb3;
	wire [3:0] la4;
	wire [3:0] lb4;
	wire [3:0] la5;
	wire [3:0] lb5;
	wire [3:0] la6;
	wire [3:0] lb6;
	wire [3:0] la7;
	wire [3:0] lb7;
	wire [3:0] la8;
	wire [3:0] lb8;
	wire [3:0] la9;
	wire [3:0] lb9;
	wire [3:0] la10;
	wire [3:0] lb10;
	wire [3:0] la11;
	wire [3:0] lb11;
	wire [3:0] la12;
	wire [3:0] lb12;
	wire [3:0] la13;
	wire [3:0] lb13;
	wire [3:0] la14;
	wire [3:0] lb14;
	wire [3:0] la15;
	wire [3:0] lb15;
	wire [3:0] la16;
	wire [3:0] lb16;
	wire [3:0] la17;
	wire [3:0] lb17;
	wire [3:0] la18;
	wire [3:0] lb18;
	wire [3:0] la19;
	wire [3:0] lb19;
	wire [3:0] la20;
	wire [3:0] lb20;
	wire [3:0] la21;
	wire [3:0] lb21;

	wire cin1;
	wire cin2;
	wire cin3;
	wire cin4;
	wire cin5;
	wire cin6;
	wire cin7;
	wire cin8;
	wire cin9;
	wire cin10;
	wire cin11;
	wire cin12;
	wire cin13;
	wire cin14;
	wire cin15;
	wire cin16;
	wire cin17;
	wire cin18;
	wire cin19;
	wire cin20;
	wire cin21;

	//Row 1
	wire [3:0] pin1;
	wire [3:0] pin2;
	wire [3:0] pin3;
	wire [3:0] pin4;
	wire [3:0] pin6;
	wire [3:0] pin7;
	wire [3:0] pin8;
	wire [3:0] pin10;
	wire [3:0] pin11;
	wire [3:0] pin12;
	wire [3:0] pin14;
	wire [3:0] pin15;
	wire [3:0] pin17;
	wire [3:0] pin18;
	wire [3:0] pin20;
	wire [3:0] pin21;
	
	
	
	wire [3:0] gin1;
	wire [3:0] gin2;
	wire [3:0] gin3;
	wire [3:0] gin4;
	wire [3:0] gin6;
	wire [3:0] gin7;
	wire [3:0] gin8;
	wire [3:0] gin10;
	wire [3:0] gin11;
	wire [3:0] gin12;
	wire [3:0] gin14;
	wire [3:0] gin15;
	wire [3:0] gin17;
	wire [3:0] gin18;
	wire [3:0] gin20;
	wire [3:0] gin21;
	
	
	// Carry LookAheads//
	//Row 1
	
	lookAheadLogic row1(cout1[2:0], gout1, pout1, pin1[3:0], gin1[3:0], cin1);
	lookAheadLogic row2(cout2[2:0], gout2, pout2, pin2[3:0], gin2[3:0], cin2);
	lookAheadLogic row3(cout3[2:0], gout3, pout3, pin3[3:0], gin3[3:0], cin3);
	lookAheadLogic row4(cout4[2:0], gout4, pout4, pin4[3:0], gin4[3:0], cin4);
	lookAheadLogic row5(cout5[2:0], gout5, pout5, la5[3:0], lb5[3:0], cin5); // gout5 is carry from row1
	pgGen pgRow1(pin1[3:0],gin1[3:0],la1,lb1);	
	pgGen pgRow2(pin2[3:0],gin2[3:0],la2,lb2);
	pgGen pgRow3(pin3[3:0],gin3[3:0],la3,lb3);
	pgGen pgRow4(pin4[3:0],gin4[3:0],la4,lb4);


	assign la1= {P_0_4,P_0_3,P_0_2,P_0_1};
	assign lb1= {P_1_3,P_1_2,P_1_1,P_1_0};
	assign cin1=0;
	assign la2= {P_0_8,P_0_7,P_0_6,P_0_5};
	assign lb2= {P_1_7,P_1_6,P_1_5,P_1_4};
	assign cin2=cout5[0];
	assign la3= {P_0_12,P_0_11,P_0_10,P_0_9};
	assign lb3= {P_1_11,P_1_10,P_1_9,P_1_8};
	assign cin3=cout5[1];
	assign la4= {2'b11,P_0_14,P_0_13};
	assign lb4= {2'b0,P_1_13,P_1_12};
	assign cin4=cout5[2];
	
	assign la5= {pout4,pout3,pout2,pout1};
	assign lb5= {gout4,gout3,gout2,gout1};
	assign cin5=0;
	
	
	
	
	
	//Row 2
	
	lookAheadLogic row6(cout6[2:0], gout6, pout6, pin6[3:0], gin6[3:0], cin6);
	lookAheadLogic row7(cout7[2:0], gout7, pout7, pin7[3:0], gin7[3:0], cin7);
	lookAheadLogic row8(cout8[2:0], gout8, pout8, pin8[3:0], gin8[3:0], cin8);
	lookAheadLogic row9(cout9[2:0], gout9, pout9, la9[3:0], lb9[3:0], cin9);// gout9 is carry from row2
	pgGen pgRow6(pin6[3:0],gin6[3:0],la6,lb6);	
	pgGen pgRow7(pin7[3:0],gin7[3:0],la7,lb7);
	pgGen pgRow8(pin8[3:0],gin8[3:0],la8,lb8);
	assign la6= {P_2_4,P_2_3,P_2_2,P_2_1};
	assign lb6= {P_3_3,P_3_2,P_3_1,P_3_0};
	assign cin6=0;
	assign la7= {P_2_8,P_2_7,P_2_6,P_2_5};
	assign lb7= {P_3_7,P_3_6,P_3_5,P_3_4};
	assign cin7=cout9[0];
	assign la8= {P_2_12,P_2_11,P_2_10,P_2_9};
	assign lb8= {P_3_11,P_3_10,P_3_9,P_3_8};
	assign cin8=cout9[1];
	
	
	assign la9= {1'b1,pout8,pout7,pout6};
	assign lb9= {1'b0,gout8,gout7,gout6};
	assign cin9=0;
	
	//Row 3
	lookAheadLogic row10(cout10[2:0], gout10, pout10, pin10[3:0], gin10[3:0], cin10);
	lookAheadLogic row11(cout11[2:0], gout11, pout11, pin11[3:0], gin11[3:0], cin11);
	lookAheadLogic row12(cout12[2:0], gout12, pout12, pin12[3:0], gin12[3:0], cin12);
	lookAheadLogic row13(cout13[2:0], gout13, pout13, la13[3:0], lb13[3:0], cin13);// gout13 is carry from row3
	pgGen pgRow10(pin10[3:0],gin10[3:0],la10,lb10);	
	pgGen pgRow11(pin11[3:0],gin11[3:0],la11,lb11);
	pgGen pgRow12(pin12[3:0],gin12[3:0],la12,lb12);
	assign la10= {P_4_4,P_4_3,P_4_2,P_4_1};
	assign lb10= {P_5_3,P_5_2,P_5_1,P_5_0};
	assign cin10=0;
	assign la11= {P_4_8,P_4_7,P_4_6,P_4_5};
	assign lb11= {P_3_7,P_3_6,P_3_5,P_3_4};
	assign cin11=cout13[0];
	assign la12= {2'b11,P_4_10,P_4_9};
	assign lb12= {2'b0,P_5_9,P_5_8};
	assign cin12=cout13[1];
	
	
	assign la13= {1'b1,pout12,pout11,pout10};
	assign lb13= {1'b0,gout12,gout11,gout10};
	assign cin13=0;
	
	//Row 4
	lookAheadLogic row14(cout14[2:0], gout14, pout14, pin14[3:0], gin14[3:0], cin14);
	lookAheadLogic row15(cout15[2:0], gout15, pout15, pin15[3:0], gin15[3:0], cin15);
	lookAheadLogic row16(cout16[2:0], gout16, pout16, la16[3:0], lb16[3:0], cin16); // gout16 is carry from row4
	pgGen pgRow14(pin14[3:0],gin14[3:0],la14,lb14);	
	pgGen pgRow15(pin15[3:0],gin15[3:0],la15,lb15);
	 
	assign la14= {P_6_4,P_6_3,P_6_2,P_6_1};
	assign lb14= {P_7_3,P_7_2,P_7_1,P_7_0};
	assign cin14=0;
	assign la15= {P_6_8,P_6_7,P_6_6,P_6_5};
	assign lb15= {P_7_7,P_7_6,P_7_5,P_7_4};
	assign cin15=cout16[0];
	
	
	
	assign la16= {2'b11,pout15,pout14};
	assign lb16= {2'b0,gout15,gout14};
	assign cin16=0;
	
	//Row 5
	lookAheadLogic row17(cout17[2:0], gout17, pout17, pin17[3:0], gin17[3:0], cin17);
	lookAheadLogic row18(cout18[2:0], gout18, pout18, pin18[3:0], gin18[3:0], cin18);
	lookAheadLogic row19(cout19[2:0], gout19, pout19, la19[3:0], lb19[3:0], cin19); // gout19 is carry from row5
	pgGen pgRow17(pin17[3:0],gin17[3:0],la17,lb17);	
	pgGen pgRow18(pin18[3:0],gin18[3:0],la18,lb18);
	 
	assign la17= {P_8_4,P_8_3,P_8_2,P_8_1};
	assign lb17= {P_9_3,P_9_2,P_9_1,P_9_0};
	assign cin17=0;
	assign la18= {2'b11,P_8_6,P_8_5};
	assign lb18= {2'b0,P_9_5,P_9_4};
	assign cin18=cout19[0];
	
	
	
	assign la19= {2'b11,pout18,pout17};
	assign lb19= {2'b0,gout18,gout17};
	assign cin19=0;
	
	//Row 6
	lookAheadLogic row20(cout20[2:0], gout20, pout20, pin20[3:0], gin20[3:0], cin20);// gout20 is carry from Row6
	pgGen pgRow20(pin20[3:0],gin20[3:0],la20,lb20);
	assign la20= {P_10_4,P_10_3,P_10_2,P_10_1};
	assign lb20= {P_11_3,P_11_2,P_11_1,P_11_0};
	assign cin20=0;
	
	//Row 7
	lookAheadLogic row21(cout21[2:0], gout21, pout21, pin21[3:0], gin21[3:0], cin21);// gout21 is carry from Row6
	pgGen pgRow21(pin21[3:0],gin21[3:0],la21,lb21);
	assign la21= {P_12_4,P_12_3,P_12_2,P_12_1};
	assign lb21= {P_13_3,P_13_2,P_13_1,P_13_0};
	assign cin21=0;


















/************************** Height - 0 ********************************/ 
//	wire S_0_0_13;
//	wire C_0_0_13;
//	halfAdder HA_0_0_13(S_0_0_13, C_0_0_13, P_0_13, P_1_12);
//	wire S_0_0_14;
//	wire C_0_0_14;
//	fullAdder FA_0_0_14(S_0_0_14, C_0_0_14, P_0_14,  P_1_13, P_2_12);
//	wire S_0_3_14;
//	wire C_0_3_14;
//	halfAdder HA_0_3_14(S_0_3_14, C_0_3_14, P_3_11, P_4_10);
	wire S_0_0_15;
	wire C_0_0_15;
	fullAdder FA_0_0_15(S_0_0_15, C_0_0_15, P_0_15,  P_1_14, P_2_13);
	wire S_0_3_15;
	wire C_0_3_15;
	fullAdder FA_0_3_15(S_0_3_15, C_0_3_15, P_3_12,  P_4_11, P_5_10);
	wire S_0_6_15;
	wire C_0_6_15;
	halfAdder HA_0_6_15(S_0_6_15, C_0_6_15, P_6_9, P_7_8);
	wire S_0_1_16;
	wire C_0_1_16;
	fullAdder FA_0_1_16(S_0_1_16, C_0_1_16, P_1_15,  P_2_14, P_3_13);
	wire S_0_4_16;
	wire C_0_4_16;
	fullAdder FA_0_4_16(S_0_4_16, C_0_4_16, P_4_12,  P_5_11, P_6_10);
	wire S_0_7_16;
	wire C_0_7_16;
	halfAdder HA_0_7_16(S_0_7_16, C_0_7_16, P_7_9, P_8_8);
	wire S_0_2_17;
	wire C_0_2_17;
	fullAdder FA_0_2_17(S_0_2_17, C_0_2_17, P_2_15,  P_3_14, P_4_13);
	wire S_0_5_17;
	wire C_0_5_17;
	fullAdder FA_0_5_17(S_0_5_17, C_0_5_17, P_5_12,  P_6_11, P_7_10);
	wire S_0_3_18;
	wire C_0_3_18;
	fullAdder FA_0_3_18(S_0_3_18, C_0_3_18, P_3_15,  P_4_14, P_5_13);
 /************************** Height - 1 ********************************/ 
//	wire S_1_0_9;
//	wire C_1_0_9;
//	halfAdder HA_1_0_9(S_1_0_9, C_1_0_9, P_0_9, P_1_8);
//	wire S_1_0_10;
//	wire C_1_0_10;
//	fullAdder FA_1_0_10(S_1_0_10, C_1_0_10, P_0_10,  P_1_9, P_2_8);
//	wire S_1_3_10;
//	wire C_1_3_10;
//	halfAdder HA_1_3_10(S_1_3_10, C_1_3_10, P_3_7, P_4_6);
//	wire S_1_0_11;
//	wire C_1_0_11;
//	fullAdder FA_1_0_11(S_1_0_11, C_1_0_11, P_0_11,  P_1_10, P_2_9);
//	wire S_1_3_11;
//	wire C_1_3_11;
//	fullAdder FA_1_3_11(S_1_3_11, C_1_3_11, P_3_8,  P_4_7, P_5_6);
//	wire S_1_6_11;
//	wire C_1_6_11;
//	halfAdder HA_1_6_11(S_1_6_11, C_1_6_11, P_6_5, P_7_4);
//	wire S_1_0_12;
//	wire C_1_0_12;
//	fullAdder FA_1_0_12(S_1_0_12, C_1_0_12, P_0_12,  P_1_11, P_2_10);
//	wire S_1_3_12;
//	wire C_1_3_12;
//	fullAdder FA_1_3_12(S_1_3_12, C_1_3_12, P_3_9,  P_4_8, P_5_7);
//	wire S_1_6_12;
//	wire C_1_6_12;
//	fullAdder FA_1_6_12(S_1_6_12, C_1_6_12, P_6_6,  P_7_5, P_8_4);
//	wire S_1_9_12;
//	wire C_1_9_12;
//	halfAdder HA_1_9_12(S_1_9_12, C_1_9_12, P_9_3, P_10_2);
//	wire S_1_0_13;
//	wire C_1_0_13;
//	fullAdder FA_1_0_13(S_1_0_13, C_1_0_13, S_0_0_13,  P_2_11, P_3_10);
//	wire S_1_3_13;
//	wire C_1_3_13;
//	fullAdder FA_1_3_13(S_1_3_13, C_1_3_13, P_4_9,  P_5_8, P_6_7);
//	wire S_1_6_13;
//	wire C_1_6_13;
//	fullAdder FA_1_6_13(S_1_6_13, C_1_6_13, P_7_6,  P_8_5, P_9_4);
//	wire S_1_9_13;
//	wire C_1_9_13;
//	fullAdder FA_1_9_13(S_1_9_13, C_1_9_13, P_10_3,  P_11_2, P_12_1);
//	wire S_1_0_14;
//	wire C_1_0_14;
//	fullAdder FA_1_0_14(S_1_0_14, C_1_0_14, C_0_0_13,  S_0_0_14, S_0_3_14);
//	wire S_1_3_14;
//	wire C_1_3_14;
//	fullAdder FA_1_3_14(S_1_3_14, C_1_3_14, P_5_9,  P_6_8, P_7_7);
//	wire S_1_6_14;
//	wire C_1_6_14;
//	fullAdder FA_1_6_14(S_1_6_14, C_1_6_14, P_8_6,  P_9_5, P_10_4);
//	wire S_1_9_14;
//	wire C_1_9_14;
//	fullAdder FA_1_9_14(S_1_9_14, C_1_9_14, P_11_3,  P_12_2, P_13_1);
	wire S_1_0_15;
	wire C_1_0_15;
	fullAdder FA_1_0_15(S_1_0_15, C_1_0_15, gout9,  gout5, S_0_0_15);	//gout5 replaces C_0_3_14 , gout9 replaces C_0_0_14
	wire S_1_3_15;
	wire C_1_3_15;
	fullAdder FA_1_3_15(S_1_3_15, C_1_3_15, S_0_3_15,  S_0_6_15, P_8_7);
	wire S_1_6_15;
	wire C_1_6_15;
	fullAdder FA_1_6_15(S_1_6_15, C_1_6_15, P_9_6,  P_10_5, P_11_4);
	wire S_1_9_15;
	wire C_1_9_15;
	fullAdder FA_1_9_15(S_1_9_15, C_1_9_15, P_12_3,  P_13_2, P_14_1);
	wire S_1_0_16;
	wire C_1_0_16;
	fullAdder FA_1_0_16(S_1_0_16, C_1_0_16, C_0_0_15,  C_0_3_15, C_0_6_15);
	wire S_1_3_16;
	wire C_1_3_16;
	fullAdder FA_1_3_16(S_1_3_16, C_1_3_16, S_0_1_16,  S_0_4_16, S_0_7_16);
	wire S_1_6_16;
	wire C_1_6_16;
	fullAdder FA_1_6_16(S_1_6_16, C_1_6_16, P_9_7,  P_10_6, P_11_5);
	wire S_1_9_16;
	wire C_1_9_16;
	fullAdder FA_1_9_16(S_1_9_16, C_1_9_16, P_12_4,  P_13_3, P_14_2);
	wire S_1_0_17;
	wire C_1_0_17;
	fullAdder FA_1_0_17(S_1_0_17, C_1_0_17, C_0_1_16,  C_0_4_16, C_0_7_16);
	wire S_1_3_17;
	wire C_1_3_17;
	fullAdder FA_1_3_17(S_1_3_17, C_1_3_17, S_0_2_17,  S_0_5_17, P_8_9);
	wire S_1_6_17;
	wire C_1_6_17;
	fullAdder FA_1_6_17(S_1_6_17, C_1_6_17, P_9_8,  P_10_7, P_11_6);
	wire S_1_9_17;
	wire C_1_9_17;
	fullAdder FA_1_9_17(S_1_9_17, C_1_9_17, P_12_5,  P_13_4, P_14_3);
	wire S_1_0_18;
	wire C_1_0_18;
	fullAdder FA_1_0_18(S_1_0_18, C_1_0_18, C_0_2_17,  C_0_5_17, S_0_3_18);
	wire S_1_3_18;
	wire C_1_3_18;
	fullAdder FA_1_3_18(S_1_3_18, C_1_3_18, P_6_12,  P_7_11, P_8_10);
	wire S_1_6_18;
	wire C_1_6_18;
	fullAdder FA_1_6_18(S_1_6_18, C_1_6_18, P_9_9,  P_10_8, P_11_7);
	wire S_1_9_18;
	wire C_1_9_18;
	fullAdder FA_1_9_18(S_1_9_18, C_1_9_18, P_12_6,  P_13_5, P_14_4);
	wire S_1_0_19;
	wire C_1_0_19;
	fullAdder FA_1_0_19(S_1_0_19, C_1_0_19, P_4_15,  P_5_14, P_6_13);
	wire S_1_3_19;
	wire C_1_3_19;
	fullAdder FA_1_3_19(S_1_3_19, C_1_3_19, P_7_12,  P_8_11, P_9_10);
	wire S_1_6_19;
	wire C_1_6_19;
	fullAdder FA_1_6_19(S_1_6_19, C_1_6_19, P_10_9,  P_11_8, P_12_7);
	wire S_1_9_19;
	wire C_1_9_19;
	fullAdder FA_1_9_19(S_1_9_19, C_1_9_19, P_13_6,  P_14_5, P_15_4);
	wire S_1_0_20;
	wire C_1_0_20;
	fullAdder FA_1_0_20(S_1_0_20, C_1_0_20, P_5_15,  P_6_14, P_7_13);
	wire S_1_3_20;
	wire C_1_3_20;
	fullAdder FA_1_3_20(S_1_3_20, C_1_3_20, P_8_12,  P_9_11, P_10_10);
	wire S_1_6_20;
	wire C_1_6_20;
	fullAdder FA_1_6_20(S_1_6_20, C_1_6_20, P_11_9,  P_12_8, P_13_7);
	wire S_1_0_21;
	wire C_1_0_21;
	fullAdder FA_1_0_21(S_1_0_21, C_1_0_21, P_6_15,  P_7_14, P_8_13);
	wire S_1_3_21;
	wire C_1_3_21;
	fullAdder FA_1_3_21(S_1_3_21, C_1_3_21, P_9_12,  P_10_11, P_11_10);
	wire S_1_0_22;
	wire C_1_0_22;
	fullAdder FA_1_0_22(S_1_0_22, C_1_0_22, P_7_15,  P_8_14, P_9_13);
 /************************** Height - 2 ********************************/ 
//	wire S_2_0_6;
//	wire C_2_0_6;
//	halfAdder HA_2_0_6(S_2_0_6, C_2_0_6, P_0_6, P_1_5);
//	wire S_2_0_7;
//	wire C_2_0_7;
//	fullAdder FA_2_0_7(S_2_0_7, C_2_0_7, P_0_7,  P_1_6, P_2_5);
//	wire S_2_3_7;
//	wire C_2_3_7;
//	halfAdder HA_2_3_7(S_2_3_7, C_2_3_7, P_3_4, P_4_3);
//	wire S_2_0_8;
//	wire C_2_0_8;
//	fullAdder FA_2_0_8(S_2_0_8, C_2_0_8, P_0_8,  P_1_7, P_2_6);
//	wire S_2_3_8;
//	wire C_2_3_8;
//	fullAdder FA_2_3_8(S_2_3_8, C_2_3_8, P_3_5,  P_4_4, P_5_3);
//	wire S_2_6_8;
//	wire C_2_6_8;
//	halfAdder HA_2_6_8(S_2_6_8, C_2_6_8, P_6_2, P_7_1);
//	wire S_2_0_9;
//	wire C_2_0_9;
//	fullAdder FA_2_0_9(S_2_0_9, C_2_0_9, S_1_0_9,  P_2_7, P_3_6);
//	wire S_2_3_9;
//	wire C_2_3_9;
//	fullAdder FA_2_3_9(S_2_3_9, C_2_3_9, P_4_5,  P_5_4, P_6_3);
//	wire S_2_6_9;
//	wire C_2_6_9;
//	fullAdder FA_2_6_9(S_2_6_9, C_2_6_9, P_7_2,  P_8_1, P_9_0);
//	wire S_2_0_10;
//	wire C_2_0_10;
//	fullAdder FA_2_0_10(S_2_0_10, C_2_0_10, C_1_0_9,  S_1_0_10, S_1_3_10);
//	wire S_2_3_10;
//	wire C_2_3_10;
//	fullAdder FA_2_3_10(S_2_3_10, C_2_3_10, P_5_5,  P_6_4, P_7_3);
//	wire S_2_6_10;
//	wire C_2_6_10;
//	fullAdder FA_2_6_10(S_2_6_10, C_2_6_10, P_8_2,  P_9_1, P_10_0);
//	wire S_2_0_11;
//	wire C_2_0_11;
//	fullAdder FA_2_0_11(S_2_0_11, C_2_0_11, C_1_0_10,  C_1_3_10, S_1_0_11);
//	wire S_2_3_11;
//	wire C_2_3_11;
//	fullAdder FA_2_3_11(S_2_3_11, C_2_3_11, S_1_3_11,  S_1_6_11, P_8_3);
//	wire S_2_6_11;
//	wire C_2_6_11;
//	fullAdder FA_2_6_11(S_2_6_11, C_2_6_11, P_9_2,  P_10_1, P_11_0);
//	wire S_2_0_12;
//	wire C_2_0_12;
//	fullAdder FA_2_0_12(S_2_0_12, C_2_0_12, C_1_0_11,  C_1_3_11, C_1_6_11);
//	wire S_2_3_12;
//	wire C_2_3_12;
//	fullAdder FA_2_3_12(S_2_3_12, C_2_3_12, S_1_0_12,  S_1_3_12, S_1_6_12);
//	wire S_2_6_12;
//	wire C_2_6_12;
//	fullAdder FA_2_6_12(S_2_6_12, C_2_6_12, S_1_9_12,  P_11_1, P_12_0);
//	wire S_2_0_13;
//	wire C_2_0_13;
//	fullAdder FA_2_0_13(S_2_0_13, C_2_0_13, C_1_0_12,  C_1_3_12, C_1_6_12);
//	wire S_2_3_13;
//	wire C_2_3_13;
//	fullAdder FA_2_3_13(S_2_3_13, C_2_3_13, C_1_9_12,  S_1_0_13, S_1_3_13);
//	wire S_2_6_13;
//	wire C_2_6_13;
//	fullAdder FA_2_6_13(S_2_6_13, C_2_6_13, S_1_6_13,  S_1_9_13, P_13_0);
//	wire S_2_0_14;
//	wire C_2_0_14;
//	fullAdder FA_2_0_14(S_2_0_14, C_2_0_14, C_1_0_13,  C_1_3_13, C_1_6_13);
//	wire S_2_3_14;
//	wire C_2_3_14;
//	fullAdder FA_2_3_14(S_2_3_14, C_2_3_14, C_1_9_13,  S_1_0_14, S_1_3_14);
//	wire S_2_6_14;
//	wire C_2_6_14;
//	fullAdder FA_2_6_14(S_2_6_14, C_2_6_14, S_1_6_14,  S_1_9_14, P_14_0);
	wire S_2_0_15;
	wire C_2_0_15;
	fullAdder FA_2_0_15(S_2_0_15, C_2_0_15, gout13,  gout16, gout19);	//gout13 replaces C_1_0_14, gout16 replaces C_1_3_14, gout19 replaces C_1_6_14
	wire S_2_3_15;
	wire C_2_3_15;
	fullAdder FA_2_3_15(S_2_3_15, C_2_3_15, gout20,  S_1_0_15, S_1_3_15);	//gout20 replaces C_1_9_14
	wire S_2_6_15;
	wire C_2_6_15;
	fullAdder FA_2_6_15(S_2_6_15, C_2_6_15, S_1_6_15,  S_1_9_15, P_15_0);
	wire S_2_0_16;
	wire C_2_0_16;
	fullAdder FA_2_0_16(S_2_0_16, C_2_0_16, C_1_0_15,  C_1_3_15, C_1_6_15);
	wire S_2_3_16;
	wire C_2_3_16;
	fullAdder FA_2_3_16(S_2_3_16, C_2_3_16, C_1_9_15,  S_1_0_16, S_1_3_16);
	wire S_2_6_16;
	wire C_2_6_16;
	fullAdder FA_2_6_16(S_2_6_16, C_2_6_16, S_1_6_16,  S_1_9_16, P_15_1);
	wire S_2_0_17;
	wire C_2_0_17;
	fullAdder FA_2_0_17(S_2_0_17, C_2_0_17, C_1_0_16,  C_1_3_16, C_1_6_16);
	wire S_2_3_17;
	wire C_2_3_17;
	fullAdder FA_2_3_17(S_2_3_17, C_2_3_17, C_1_9_16,  S_1_0_17, S_1_3_17);
	wire S_2_6_17;
	wire C_2_6_17;
	fullAdder FA_2_6_17(S_2_6_17, C_2_6_17, S_1_6_17,  S_1_9_17, P_15_2);
	wire S_2_0_18;
	wire C_2_0_18;
	fullAdder FA_2_0_18(S_2_0_18, C_2_0_18, C_1_0_17,  C_1_3_17, C_1_6_17);
	wire S_2_3_18;
	wire C_2_3_18;
	fullAdder FA_2_3_18(S_2_3_18, C_2_3_18, C_1_9_17,  S_1_0_18, S_1_3_18);
	wire S_2_6_18;
	wire C_2_6_18;
	fullAdder FA_2_6_18(S_2_6_18, C_2_6_18, S_1_6_18,  S_1_9_18, P_15_3);
	wire S_2_0_19;
	wire C_2_0_19;
	fullAdder FA_2_0_19(S_2_0_19, C_2_0_19, C_1_0_18,  C_1_3_18, C_1_6_18);
	wire S_2_3_19;
	wire C_2_3_19;
	fullAdder FA_2_3_19(S_2_3_19, C_2_3_19, C_1_9_18,  S_1_0_19, S_1_3_19);
	wire S_2_6_19;
	wire C_2_6_19;
	fullAdder FA_2_6_19(S_2_6_19, C_2_6_19, S_1_6_19,  S_1_9_19, C_0_3_18);
	wire S_2_0_20;
	wire C_2_0_20;
	fullAdder FA_2_0_20(S_2_0_20, C_2_0_20, C_1_0_19,  C_1_3_19, C_1_6_19);
	wire S_2_3_20;
	wire C_2_3_20;
	fullAdder FA_2_3_20(S_2_3_20, C_2_3_20, C_1_9_19,  S_1_0_20, S_1_3_20);
	wire S_2_6_20;
	wire C_2_6_20;
	fullAdder FA_2_6_20(S_2_6_20, C_2_6_20, S_1_6_20,  P_14_6, P_15_5);
	wire S_2_0_21;
	wire C_2_0_21;
	fullAdder FA_2_0_21(S_2_0_21, C_2_0_21, C_1_0_20,  C_1_3_20, C_1_6_20);
	wire S_2_3_21;
	wire C_2_3_21;
	fullAdder FA_2_3_21(S_2_3_21, C_2_3_21, S_1_0_21,  S_1_3_21, P_12_9);
	wire S_2_6_21;
	wire C_2_6_21;
	fullAdder FA_2_6_21(S_2_6_21, C_2_6_21, P_13_8,  P_14_7, P_15_6);
	wire S_2_0_22;
	wire C_2_0_22;
	fullAdder FA_2_0_22(S_2_0_22, C_2_0_22, C_1_0_21,  C_1_3_21, S_1_0_22);
	wire S_2_3_22;
	wire C_2_3_22;
	fullAdder FA_2_3_22(S_2_3_22, C_2_3_22, P_10_12,  P_11_11, P_12_10);
	wire S_2_6_22;
	wire C_2_6_22;
	fullAdder FA_2_6_22(S_2_6_22, C_2_6_22, P_13_9,  P_14_8, P_15_7);
	wire S_2_0_23;
	wire C_2_0_23;
	fullAdder FA_2_0_23(S_2_0_23, C_2_0_23, P_8_15,  P_9_14, P_10_13);
	wire S_2_3_23;
	wire C_2_3_23;
	fullAdder FA_2_3_23(S_2_3_23, C_2_3_23, P_11_12,  P_12_11, P_13_10);
	wire S_2_6_23;
	wire C_2_6_23;
	fullAdder FA_2_6_23(S_2_6_23, C_2_6_23, P_14_9,  P_15_8, C_1_0_22);
	wire S_2_0_24;
	wire C_2_0_24;
	fullAdder FA_2_0_24(S_2_0_24, C_2_0_24, P_9_15,  P_10_14, P_11_13);
	wire S_2_3_24;
	wire C_2_3_24;
	fullAdder FA_2_3_24(S_2_3_24, C_2_3_24, P_12_12,  P_13_11, P_14_10);
	wire S_2_0_25;
	wire C_2_0_25;
	fullAdder FA_2_0_25(S_2_0_25, C_2_0_25, P_10_15,  P_11_14, P_12_13);
 /************************** Height - 3 ********************************/ 
//	wire S_3_0_4;
//	wire C_3_0_4;
//	halfAdder HA_3_0_4(S_3_0_4, C_3_0_4, P_0_4, P_1_3);
//	wire S_3_0_5;
//	wire C_3_0_5;
//	fullAdder FA_3_0_5(S_3_0_5, C_3_0_5, P_0_5,  P_1_4, P_2_3);
//	wire S_3_3_5;
//	wire C_3_3_5;
//	halfAdder HA_3_3_5(S_3_3_5, C_3_3_5, P_3_2, P_4_1);
//	wire S_3_0_6;
//	wire C_3_0_6;
//	fullAdder FA_3_0_6(S_3_0_6, C_3_0_6, S_2_0_6,  P_2_4, P_3_3);
//	wire S_3_3_6;
//	wire C_3_3_6;
//	fullAdder FA_3_3_6(S_3_3_6, C_3_3_6, P_4_2,  P_5_1, P_6_0);
//	wire S_3_0_7;
//	wire C_3_0_7;
//	fullAdder FA_3_0_7(S_3_0_7, C_3_0_7, C_2_0_6,  S_2_0_7, S_2_3_7);
//	wire S_3_3_7;
//	wire C_3_3_7;
//	fullAdder FA_3_3_7(S_3_3_7, C_3_3_7, P_5_2,  P_6_1, P_7_0);
//	wire S_3_0_8;
//	wire C_3_0_8;
//	fullAdder FA_3_0_8(S_3_0_8, C_3_0_8, C_2_0_7,  C_2_3_7, S_2_0_8);
//	wire S_3_3_8;
//	wire C_3_3_8;
//	fullAdder FA_3_3_8(S_3_3_8, C_3_3_8, S_2_3_8,  S_2_6_8, P_8_0);
//	wire S_3_0_9;
//	wire C_3_0_9;
//	fullAdder FA_3_0_9(S_3_0_9, C_3_0_9, C_2_0_8,  C_2_3_8, C_2_6_8);
//	wire S_3_3_9;
//	wire C_3_3_9;
//	fullAdder FA_3_3_9(S_3_3_9, C_3_3_9, S_2_0_9,  S_2_3_9, S_2_6_9);
//	wire S_3_0_10;
//	wire C_3_0_10;
//	fullAdder FA_3_0_10(S_3_0_10, C_3_0_10, C_2_0_9,  C_2_3_9, C_2_6_9);
//	wire S_3_3_10;
//	wire C_3_3_10;
//	fullAdder FA_3_3_10(S_3_3_10, C_3_3_10, S_2_0_10,  S_2_3_10, S_2_6_10);
//	wire S_3_0_11;
//	wire C_3_0_11;
//	fullAdder FA_3_0_11(S_3_0_11, C_3_0_11, C_2_0_10,  C_2_3_10, C_2_6_10);
//	wire S_3_3_11;
//	wire C_3_3_11;
//	fullAdder FA_3_3_11(S_3_3_11, C_3_3_11, S_2_0_11,  S_2_3_11, S_2_6_11);
//	wire S_3_0_12;
//	wire C_3_0_12;
//	fullAdder FA_3_0_12(S_3_0_12, C_3_0_12, C_2_0_11,  C_2_3_11, C_2_6_11);
//	wire S_3_3_12;
//	wire C_3_3_12;
//	fullAdder FA_3_3_12(S_3_3_12, C_3_3_12, S_2_0_12,  S_2_3_12, S_2_6_12);
//	wire S_3_0_13;
//	wire C_3_0_13;
//	fullAdder FA_3_0_13(S_3_0_13, C_3_0_13, C_2_0_12,  C_2_3_12, C_2_6_12);
//	wire S_3_3_13;
//	wire C_3_3_13;
//	fullAdder FA_3_3_13(S_3_3_13, C_3_3_13, S_2_0_13,  S_2_3_13, S_2_6_13);
//	wire S_3_0_14;
//	wire C_3_0_14;
//	fullAdder FA_3_0_14(S_3_0_14, C_3_0_14, C_2_0_13,  C_2_3_13, C_2_6_13);
//	wire S_3_3_14;
//	wire C_3_3_14;
//	fullAdder FA_3_3_14(S_3_3_14, C_3_3_14, S_2_0_14,  S_2_3_14, S_2_6_14);
	wire S_3_0_15;
	wire C_3_0_15;
//	fullAdder FA_3_0_15(S_3_0_15, C_3_0_15, gout21,  C_2_3_14, C_2_6_14);		//gout21 replaces C_2_0_14
	assign S_3_0_15		= gout21;
	assign C_3_0_15		= 1'b0;
	wire S_3_3_15;
	wire C_3_3_15;
	fullAdder FA_3_3_15(S_3_3_15, C_3_3_15, S_2_0_15,  S_2_3_15, S_2_6_15);
	wire S_3_0_16;
	wire C_3_0_16;
	fullAdder FA_3_0_16(S_3_0_16, C_3_0_16, C_2_0_15,  C_2_3_15, C_2_6_15);
	wire S_3_3_16;
	wire C_3_3_16;
	fullAdder FA_3_3_16(S_3_3_16, C_3_3_16, S_2_0_16,  S_2_3_16, S_2_6_16);
	wire S_3_0_17;
	wire C_3_0_17;
	fullAdder FA_3_0_17(S_3_0_17, C_3_0_17, C_2_0_16,  C_2_3_16, C_2_6_16);
	wire S_3_3_17;
	wire C_3_3_17;
	fullAdder FA_3_3_17(S_3_3_17, C_3_3_17, S_2_0_17,  S_2_3_17, S_2_6_17);
	wire S_3_0_18;
	wire C_3_0_18;
	fullAdder FA_3_0_18(S_3_0_18, C_3_0_18, C_2_0_17,  C_2_3_17, C_2_6_17);
	wire S_3_3_18;
	wire C_3_3_18;
	fullAdder FA_3_3_18(S_3_3_18, C_3_3_18, S_2_0_18,  S_2_3_18, S_2_6_18);
	wire S_3_0_19;
	wire C_3_0_19;
	fullAdder FA_3_0_19(S_3_0_19, C_3_0_19, C_2_0_18,  C_2_3_18, C_2_6_18);
	wire S_3_3_19;
	wire C_3_3_19;
	fullAdder FA_3_3_19(S_3_3_19, C_3_3_19, S_2_0_19,  S_2_3_19, S_2_6_19);
	wire S_3_0_20;
	wire C_3_0_20;
	fullAdder FA_3_0_20(S_3_0_20, C_3_0_20, C_2_0_19,  C_2_3_19, C_2_6_19);
	wire S_3_3_20;
	wire C_3_3_20;
	fullAdder FA_3_3_20(S_3_3_20, C_3_3_20, S_2_0_20,  S_2_3_20, S_2_6_20);
	wire S_3_0_21;
	wire C_3_0_21;
	fullAdder FA_3_0_21(S_3_0_21, C_3_0_21, C_2_0_20,  C_2_3_20, C_2_6_20);
	wire S_3_3_21;
	wire C_3_3_21;
	fullAdder FA_3_3_21(S_3_3_21, C_3_3_21, S_2_0_21,  S_2_3_21, S_2_6_21);
	wire S_3_0_22;
	wire C_3_0_22;
	fullAdder FA_3_0_22(S_3_0_22, C_3_0_22, C_2_0_21,  C_2_3_21, C_2_6_21);
	wire S_3_3_22;
	wire C_3_3_22;
	fullAdder FA_3_3_22(S_3_3_22, C_3_3_22, S_2_0_22,  S_2_3_22, S_2_6_22);
	wire S_3_0_23;
	wire C_3_0_23;
	fullAdder FA_3_0_23(S_3_0_23, C_3_0_23, C_2_0_22,  C_2_3_22, C_2_6_22);
	wire S_3_3_23;
	wire C_3_3_23;
	fullAdder FA_3_3_23(S_3_3_23, C_3_3_23, S_2_0_23,  S_2_3_23, S_2_6_23);
	wire S_3_0_24;
	wire C_3_0_24;
	fullAdder FA_3_0_24(S_3_0_24, C_3_0_24, C_2_0_23,  C_2_3_23, C_2_6_23);
	wire S_3_3_24;
	wire C_3_3_24;
	fullAdder FA_3_3_24(S_3_3_24, C_3_3_24, S_2_0_24,  S_2_3_24, P_15_9);
	wire S_3_0_25;
	wire C_3_0_25;
	fullAdder FA_3_0_25(S_3_0_25, C_3_0_25, C_2_0_24,  C_2_3_24, S_2_0_25);
	wire S_3_3_25;
	wire C_3_3_25;
	fullAdder FA_3_3_25(S_3_3_25, C_3_3_25, P_13_12,  P_14_11, P_15_10);
	wire S_3_0_26;
	wire C_3_0_26;
	fullAdder FA_3_0_26(S_3_0_26, C_3_0_26, P_11_15,  P_12_14, P_13_13);
	wire S_3_3_26;
	wire C_3_3_26;
	fullAdder FA_3_3_26(S_3_3_26, C_3_3_26, P_14_12,  P_15_11, C_2_0_25);
	wire S_3_0_27;
	wire C_3_0_27;
	fullAdder FA_3_0_27(S_3_0_27, C_3_0_27, P_12_15,  P_13_14, P_14_13);
 /************************** Height - 4 ********************************/ 
//	wire S_4_0_3;
//	wire C_4_0_3;
//	halfAdder HA_4_0_3(S_4_0_3, C_4_0_3, P_0_3, P_1_2);
//	wire S_4_0_4;
//	wire C_4_0_4;
//	fullAdder FA_4_0_4(S_4_0_4, C_4_0_4, S_3_0_4,  P_2_2, P_3_1);
//	wire S_4_0_5;
//	wire C_4_0_5;
//	fullAdder FA_4_0_5(S_4_0_5, C_4_0_5, C_3_0_4,  S_3_0_5, S_3_3_5);
//	wire S_4_0_6;
//	wire C_4_0_6;
//	fullAdder FA_4_0_6(S_4_0_6, C_4_0_6, C_3_0_5,  C_3_3_5, S_3_0_6);
//	wire S_4_0_7;
//	wire C_4_0_7;
//	fullAdder FA_4_0_7(S_4_0_7, C_4_0_7, C_3_0_6,  C_3_3_6, S_3_0_7);
//	wire S_4_0_8;
//	wire C_4_0_8;
//	fullAdder FA_4_0_8(S_4_0_8, C_4_0_8, C_3_0_7,  C_3_3_7, S_3_0_8);
//	wire S_4_0_9;
//	wire C_4_0_9;
//	fullAdder FA_4_0_9(S_4_0_9, C_4_0_9, C_3_0_8,  C_3_3_8, S_3_0_9);
//	wire S_4_0_10;
//	wire C_4_0_10;
//	fullAdder FA_4_0_10(S_4_0_10, C_4_0_10, C_3_0_9,  C_3_3_9, S_3_0_10);
//	wire S_4_0_11;
//	wire C_4_0_11;
//	fullAdder FA_4_0_11(S_4_0_11, C_4_0_11, C_3_0_10,  C_3_3_10, S_3_0_11);
//	wire S_4_0_12;
//	wire C_4_0_12;
//	fullAdder FA_4_0_12(S_4_0_12, C_4_0_12, C_3_0_11,  C_3_3_11, S_3_0_12);
//	wire S_4_0_13;
//	wire C_4_0_13;
//	fullAdder FA_4_0_13(S_4_0_13, C_4_0_13, C_3_0_12,  C_3_3_12, S_3_0_13);
//	wire S_4_0_14;
//	wire C_4_0_14;
//	fullAdder FA_4_0_14(S_4_0_14, C_4_0_14, C_3_0_13,  C_3_3_13, S_3_0_14);
	wire S_4_0_15;
	wire C_4_0_15;
	assign S_4_0_15		= S_3_0_15;
	assign C_4_0_15		= 1'b0;
//	fullAdder FA_4_0_15(S_4_0_15, C_4_0_15, C_3_0_14,  1'b0, S_3_0_15);
	wire S_4_0_16;
	wire C_4_0_16;
	halfAdder HA_4_0_16(S_4_0_16, C_4_0_16, C_3_3_15, S_3_0_16);
	wire S_4_0_17;
	wire C_4_0_17;
	fullAdder FA_4_0_17(S_4_0_17, C_4_0_17, C_3_0_16,  C_3_3_16, S_3_0_17);
	wire S_4_0_18;
	wire C_4_0_18;
	fullAdder FA_4_0_18(S_4_0_18, C_4_0_18, C_3_0_17,  C_3_3_17, S_3_0_18);
	wire S_4_0_19;
	wire C_4_0_19;
	fullAdder FA_4_0_19(S_4_0_19, C_4_0_19, C_3_0_18,  C_3_3_18, S_3_0_19);
	wire S_4_0_20;
	wire C_4_0_20;
	fullAdder FA_4_0_20(S_4_0_20, C_4_0_20, C_3_0_19,  C_3_3_19, S_3_0_20);
	wire S_4_0_21;
	wire C_4_0_21;
	fullAdder FA_4_0_21(S_4_0_21, C_4_0_21, C_3_0_20,  C_3_3_20, S_3_0_21);
	wire S_4_0_22;
	wire C_4_0_22;
	fullAdder FA_4_0_22(S_4_0_22, C_4_0_22, C_3_0_21,  C_3_3_21, S_3_0_22);
	wire S_4_0_23;
	wire C_4_0_23;
	fullAdder FA_4_0_23(S_4_0_23, C_4_0_23, C_3_0_22,  C_3_3_22, S_3_0_23);
	wire S_4_0_24;
	wire C_4_0_24;
	fullAdder FA_4_0_24(S_4_0_24, C_4_0_24, C_3_0_23,  C_3_3_23, S_3_0_24);
	wire S_4_0_25;
	wire C_4_0_25;
	fullAdder FA_4_0_25(S_4_0_25, C_4_0_25, C_3_0_24,  C_3_3_24, S_3_0_25);
	wire S_4_0_26;
	wire C_4_0_26;
	fullAdder FA_4_0_26(S_4_0_26, C_4_0_26, C_3_0_25,  C_3_3_25, S_3_0_26);
	wire S_4_0_27;
	wire C_4_0_27;
	fullAdder FA_4_0_27(S_4_0_27, C_4_0_27, C_3_0_26,  C_3_3_26, S_3_0_27);
	wire S_4_0_28;
	wire C_4_0_28;
	fullAdder FA_4_0_28(S_4_0_28, C_4_0_28, P_13_15,  P_14_14, P_15_13);
 /************************** Height - 5 ********************************/ 
//	wire S_5_0_2;
//	wire C_5_0_2;
//	halfAdder HA_5_0_2(S_5_0_2, C_5_0_2, P_0_2, P_1_1);
//	wire S_5_0_3;
//	wire C_5_0_3;
//	fullAdder FA_5_0_3(S_5_0_3, C_5_0_3, S_4_0_3,  P_2_1, P_3_0);
//	wire S_5_0_4;
//	wire C_5_0_4;
//	fullAdder FA_5_0_4(S_5_0_4, C_5_0_4, C_4_0_3,  S_4_0_4, P_4_0);
//	wire S_5_0_5;
//	wire C_5_0_5;
//	fullAdder FA_5_0_5(S_5_0_5, C_5_0_5, C_4_0_4,  S_4_0_5, P_5_0);
//	wire S_5_0_6;
//	wire C_5_0_6;
//	fullAdder FA_5_0_6(S_5_0_6, C_5_0_6, C_4_0_5,  S_4_0_6, S_3_3_6);
//	wire S_5_0_7;
//	wire C_5_0_7;
//	fullAdder FA_5_0_7(S_5_0_7, C_5_0_7, C_4_0_6,  S_4_0_7, S_3_3_7);
//	wire S_5_0_8;
//	wire C_5_0_8;
//	fullAdder FA_5_0_8(S_5_0_8, C_5_0_8, C_4_0_7,  S_4_0_8, S_3_3_8);
//	wire S_5_0_9;
//	wire C_5_0_9;
//	fullAdder FA_5_0_9(S_5_0_9, C_5_0_9, C_4_0_8,  S_4_0_9, S_3_3_9);
//	wire S_5_0_10;
//	wire C_5_0_10;
//	fullAdder FA_5_0_10(S_5_0_10, C_5_0_10, C_4_0_9,  S_4_0_10, S_3_3_10);
//	wire S_5_0_11;
//	wire C_5_0_11;
//	fullAdder FA_5_0_11(S_5_0_11, C_5_0_11, C_4_0_10,  S_4_0_11, S_3_3_11);
//	wire S_5_0_12;
//	wire C_5_0_12;
//	fullAdder FA_5_0_12(S_5_0_12, C_5_0_12, C_4_0_11,  S_4_0_12, S_3_3_12);
//	wire S_5_0_13;
//	wire C_5_0_13;
//	fullAdder FA_5_0_13(S_5_0_13, C_5_0_13, C_4_0_12,  S_4_0_13, S_3_3_13);
//	wire S_5_0_14;
//	wire C_5_0_14;
//	fullAdder FA_5_0_14(S_5_0_14, C_5_0_14, C_4_0_13,  S_4_0_14, S_3_3_14);
	wire S_5_0_15;
	wire C_5_0_15;
	halfAdder HA_5_0_15(S_5_0_15, C_5_0_15, S_4_0_15, S_3_3_15);
	wire S_5_0_16;
	wire C_5_0_16;
	fullAdder FA_5_0_16(S_5_0_16, C_5_0_16, C_4_0_15,  S_4_0_16, S_3_3_16);
	wire S_5_0_17;
	wire C_5_0_17;
	fullAdder FA_5_0_17(S_5_0_17, C_5_0_17, C_4_0_16,  S_4_0_17, S_3_3_17);
	wire S_5_0_18;
	wire C_5_0_18;
	fullAdder FA_5_0_18(S_5_0_18, C_5_0_18, C_4_0_17,  S_4_0_18, S_3_3_18);
	wire S_5_0_19;
	wire C_5_0_19;
	fullAdder FA_5_0_19(S_5_0_19, C_5_0_19, C_4_0_18,  S_4_0_19, S_3_3_19);
	wire S_5_0_20;
	wire C_5_0_20;
	fullAdder FA_5_0_20(S_5_0_20, C_5_0_20, C_4_0_19,  S_4_0_20, S_3_3_20);
	wire S_5_0_21;
	wire C_5_0_21;
	fullAdder FA_5_0_21(S_5_0_21, C_5_0_21, C_4_0_20,  S_4_0_21, S_3_3_21);
	wire S_5_0_22;
	wire C_5_0_22;
	fullAdder FA_5_0_22(S_5_0_22, C_5_0_22, C_4_0_21,  S_4_0_22, S_3_3_22);
	wire S_5_0_23;
	wire C_5_0_23;
	fullAdder FA_5_0_23(S_5_0_23, C_5_0_23, C_4_0_22,  S_4_0_23, S_3_3_23);
	wire S_5_0_24;
	wire C_5_0_24;
	fullAdder FA_5_0_24(S_5_0_24, C_5_0_24, C_4_0_23,  S_4_0_24, S_3_3_24);
	wire S_5_0_25;
	wire C_5_0_25;
	fullAdder FA_5_0_25(S_5_0_25, C_5_0_25, C_4_0_24,  S_4_0_25, S_3_3_25);
	wire S_5_0_26;
	wire C_5_0_26;
	fullAdder FA_5_0_26(S_5_0_26, C_5_0_26, C_4_0_25,  S_4_0_26, S_3_3_26);
	wire S_5_0_27;
	wire C_5_0_27;
	fullAdder FA_5_0_27(S_5_0_27, C_5_0_27, C_4_0_26,  S_4_0_27, P_15_12);
	wire S_5_0_28;
	wire C_5_0_28;
	fullAdder FA_5_0_28(S_5_0_28, C_5_0_28, C_4_0_27,  S_4_0_28, C_3_0_27);
	wire S_5_0_29;
	wire C_5_0_29;
	fullAdder FA_5_0_29(S_5_0_29, C_5_0_29, P_14_15,  P_15_14, C_4_0_28);
	
	
	wire [15:0] in1 = {P_15_15,S_5_0_29,S_5_0_28,S_5_0_27,S_5_0_26,S_5_0_25,S_5_0_24,S_5_0_23,S_5_0_22,S_5_0_21,S_5_0_20,S_5_0_19,S_5_0_18,S_5_0_17,S_5_0_16};
	wire [15:0] in2 = {C_5_0_29,C_5_0_28,C_5_0_27,C_5_0_26,C_5_0_25,C_5_0_24,C_5_0_23,C_5_0_22,C_5_0_21,C_5_0_20,C_5_0_19,C_5_0_18,C_5_0_17,C_5_0_16,C_5_0_15};
	
	
	assign out= in1+in2;
	assign out_end = S_5_0_15;
	
endmodule
	

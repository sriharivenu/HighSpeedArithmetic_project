module dadda8_orig(out, a, b);

	input [7:0] a;
	input [7:0] b;
	output [15:0] out;


 /************************** AND gate DOT PRODUCT matrix ********************************/ 
	wire P_0_0;
	and A_0_0(P_0_0, a[0], b[0]);
	wire P_0_1;
	and A_0_1(P_0_1, a[0], b[1]);
	wire P_0_2;
	and A_0_2(P_0_2, a[0], b[2]);
	wire P_0_3;
	and A_0_3(P_0_3, a[0], b[3]);
	wire P_0_4;
	and A_0_4(P_0_4, a[0], b[4]);
	wire P_0_5;
	and A_0_5(P_0_5, a[0], b[5]);
	wire P_0_6;
	and A_0_6(P_0_6, a[0], b[6]);
	wire P_0_7;
	and A_0_7(P_0_7, a[0], b[7]);
	wire P_1_0;
	and A_1_0(P_1_0, a[1], b[0]);
	wire P_1_1;
	and A_1_1(P_1_1, a[1], b[1]);
	wire P_1_2;
	and A_1_2(P_1_2, a[1], b[2]);
	wire P_1_3;
	and A_1_3(P_1_3, a[1], b[3]);
	wire P_1_4;
	and A_1_4(P_1_4, a[1], b[4]);
	wire P_1_5;
	and A_1_5(P_1_5, a[1], b[5]);
	wire P_1_6;
	and A_1_6(P_1_6, a[1], b[6]);
	wire P_1_7;
	and A_1_7(P_1_7, a[1], b[7]);
	wire P_2_0;
	and A_2_0(P_2_0, a[2], b[0]);
	wire P_2_1;
	and A_2_1(P_2_1, a[2], b[1]);
	wire P_2_2;
	and A_2_2(P_2_2, a[2], b[2]);
	wire P_2_3;
	and A_2_3(P_2_3, a[2], b[3]);
	wire P_2_4;
	and A_2_4(P_2_4, a[2], b[4]);
	wire P_2_5;
	and A_2_5(P_2_5, a[2], b[5]);
	wire P_2_6;
	and A_2_6(P_2_6, a[2], b[6]);
	wire P_2_7;
	and A_2_7(P_2_7, a[2], b[7]);
	wire P_3_0;
	and A_3_0(P_3_0, a[3], b[0]);
	wire P_3_1;
	and A_3_1(P_3_1, a[3], b[1]);
	wire P_3_2;
	and A_3_2(P_3_2, a[3], b[2]);
	wire P_3_3;
	and A_3_3(P_3_3, a[3], b[3]);
	wire P_3_4;
	and A_3_4(P_3_4, a[3], b[4]);
	wire P_3_5;
	and A_3_5(P_3_5, a[3], b[5]);
	wire P_3_6;
	and A_3_6(P_3_6, a[3], b[6]);
	wire P_3_7;
	and A_3_7(P_3_7, a[3], b[7]);
	wire P_4_0;
	and A_4_0(P_4_0, a[4], b[0]);
	wire P_4_1;
	and A_4_1(P_4_1, a[4], b[1]);
	wire P_4_2;
	and A_4_2(P_4_2, a[4], b[2]);
	wire P_4_3;
	and A_4_3(P_4_3, a[4], b[3]);
	wire P_4_4;
	and A_4_4(P_4_4, a[4], b[4]);
	wire P_4_5;
	and A_4_5(P_4_5, a[4], b[5]);
	wire P_4_6;
	and A_4_6(P_4_6, a[4], b[6]);
	wire P_4_7;
	and A_4_7(P_4_7, a[4], b[7]);
	wire P_5_0;
	and A_5_0(P_5_0, a[5], b[0]);
	wire P_5_1;
	and A_5_1(P_5_1, a[5], b[1]);
	wire P_5_2;
	and A_5_2(P_5_2, a[5], b[2]);
	wire P_5_3;
	and A_5_3(P_5_3, a[5], b[3]);
	wire P_5_4;
	and A_5_4(P_5_4, a[5], b[4]);
	wire P_5_5;
	and A_5_5(P_5_5, a[5], b[5]);
	wire P_5_6;
	and A_5_6(P_5_6, a[5], b[6]);
	wire P_5_7;
	and A_5_7(P_5_7, a[5], b[7]);
	wire P_6_0;
	and A_6_0(P_6_0, a[6], b[0]);
	wire P_6_1;
	and A_6_1(P_6_1, a[6], b[1]);
	wire P_6_2;
	and A_6_2(P_6_2, a[6], b[2]);
	wire P_6_3;
	and A_6_3(P_6_3, a[6], b[3]);
	wire P_6_4;
	and A_6_4(P_6_4, a[6], b[4]);
	wire P_6_5;
	and A_6_5(P_6_5, a[6], b[5]);
	wire P_6_6;
	and A_6_6(P_6_6, a[6], b[6]);
	wire P_6_7;
	and A_6_7(P_6_7, a[6], b[7]);
	wire P_7_0;
	and A_7_0(P_7_0, a[7], b[0]);
	wire P_7_1;
	and A_7_1(P_7_1, a[7], b[1]);
	wire P_7_2;
	and A_7_2(P_7_2, a[7], b[2]);
	wire P_7_3;
	and A_7_3(P_7_3, a[7], b[3]);
	wire P_7_4;
	and A_7_4(P_7_4, a[7], b[4]);
	wire P_7_5;
	and A_7_5(P_7_5, a[7], b[5]);
	wire P_7_6;
	and A_7_6(P_7_6, a[7], b[6]);
	wire P_7_7;
	and A_7_7(P_7_7, a[7], b[7]);
 /************************** Height - 0 ********************************/ 
	wire S_0_0_6;
	wire C_0_0_6;
	halfAdder HA_0_0_6(S_0_0_6, C_0_0_6, P_0_6, P_1_5);
	wire S_0_0_7;
	wire C_0_0_7;
	fullAdder FA_0_0_7(S_0_0_7, C_0_0_7, P_0_7,  P_1_6, P_2_5);
	wire S_0_3_7;
	wire C_0_3_7;
	halfAdder HA_0_3_7(S_0_3_7, C_0_3_7, P_3_4, P_4_3);
	wire S_0_1_8;
	wire C_0_1_8;
	fullAdder FA_0_1_8(S_0_1_8, C_0_1_8, P_1_7,  P_2_6, P_3_5);
	wire S_0_4_8;
	wire C_0_4_8;
	halfAdder HA_0_4_8(S_0_4_8, C_0_4_8, P_4_4, P_5_3);
	wire S_0_2_9;
	wire C_0_2_9;
	fullAdder FA_0_2_9(S_0_2_9, C_0_2_9, P_2_7,  P_3_6, P_4_5);
 /************************** Height - 1 ********************************/ 
	wire S_1_0_4;
	wire C_1_0_4;
	halfAdder HA_1_0_4(S_1_0_4, C_1_0_4, P_0_4, P_1_3);
	wire S_1_0_5;
	wire C_1_0_5;
	fullAdder FA_1_0_5(S_1_0_5, C_1_0_5, P_0_5,  P_1_4, P_2_3);
	wire S_1_3_5;
	wire C_1_3_5;
	halfAdder HA_1_3_5(S_1_3_5, C_1_3_5, P_3_2, P_4_1);
	wire S_1_0_6;
	wire C_1_0_6;
	fullAdder FA_1_0_6(S_1_0_6, C_1_0_6, S_0_0_6,  P_2_4, P_3_3);
	wire S_1_3_6;
	wire C_1_3_6;
	fullAdder FA_1_3_6(S_1_3_6, C_1_3_6, P_4_2,  P_5_1, P_6_0);
	wire S_1_0_7;
	wire C_1_0_7;
	fullAdder FA_1_0_7(S_1_0_7, C_1_0_7, C_0_0_6,  S_0_0_7, S_0_3_7);
	wire S_1_3_7;
	wire C_1_3_7;
	fullAdder FA_1_3_7(S_1_3_7, C_1_3_7, P_5_2,  P_6_1, P_7_0);
	wire S_1_0_8;
	wire C_1_0_8;
	fullAdder FA_1_0_8(S_1_0_8, C_1_0_8, C_0_0_7,  C_0_3_7, S_0_1_8);
	wire S_1_3_8;
	wire C_1_3_8;
	fullAdder FA_1_3_8(S_1_3_8, C_1_3_8, S_0_4_8,  P_6_2, P_7_1);
	wire S_1_0_9;
	wire C_1_0_9;
	fullAdder FA_1_0_9(S_1_0_9, C_1_0_9, C_0_1_8,  C_0_4_8, S_0_2_9);
	wire S_1_3_9;
	wire C_1_3_9;
	fullAdder FA_1_3_9(S_1_3_9, C_1_3_9, P_5_4,  P_6_3, P_7_2);
	wire S_1_0_10;
	wire C_1_0_10;
	fullAdder FA_1_0_10(S_1_0_10, C_1_0_10, P_3_7,  P_4_6, P_5_5);
	wire S_1_3_10;
	wire C_1_3_10;
	fullAdder FA_1_3_10(S_1_3_10, C_1_3_10, P_6_4,  P_7_3, C_0_2_9);
	wire S_1_0_11;
	wire C_1_0_11;
	fullAdder FA_1_0_11(S_1_0_11, C_1_0_11, P_4_7,  P_5_6, P_6_5);
 /************************** Height - 2 ********************************/ 
	wire S_2_0_3;
	wire C_2_0_3;
	halfAdder HA_2_0_3(S_2_0_3, C_2_0_3, P_0_3, P_1_2);
	wire S_2_0_4;
	wire C_2_0_4;
	fullAdder FA_2_0_4(S_2_0_4, C_2_0_4, S_1_0_4,  P_2_2, P_3_1);
	wire S_2_0_5;
	wire C_2_0_5;
	fullAdder FA_2_0_5(S_2_0_5, C_2_0_5, C_1_0_4,  S_1_0_5, S_1_3_5);
	wire S_2_0_6;
	wire C_2_0_6;
	fullAdder FA_2_0_6(S_2_0_6, C_2_0_6, C_1_0_5,  C_1_3_5, S_1_0_6);
	wire S_2_0_7;
	wire C_2_0_7;
	fullAdder FA_2_0_7(S_2_0_7, C_2_0_7, C_1_0_6,  C_1_3_6, S_1_0_7);
	wire S_2_0_8;
	wire C_2_0_8;
	fullAdder FA_2_0_8(S_2_0_8, C_2_0_8, C_1_0_7,  C_1_3_7, S_1_0_8);
	wire S_2_0_9;
	wire C_2_0_9;
	fullAdder FA_2_0_9(S_2_0_9, C_2_0_9, C_1_0_8,  C_1_3_8, S_1_0_9);
	wire S_2_0_10;
	wire C_2_0_10;
	fullAdder FA_2_0_10(S_2_0_10, C_2_0_10, C_1_0_9,  C_1_3_9, S_1_0_10);
	wire S_2_0_11;
	wire C_2_0_11;
	fullAdder FA_2_0_11(S_2_0_11, C_2_0_11, C_1_0_10,  C_1_3_10, S_1_0_11);
	wire S_2_0_12;
	wire C_2_0_12;
	fullAdder FA_2_0_12(S_2_0_12, C_2_0_12, P_5_7,  P_6_6, P_7_5);
 /************************** Height - 3 ********************************/ 
	wire S_3_0_2;
	wire C_3_0_2;
	halfAdder HA_3_0_2(S_3_0_2, C_3_0_2, P_0_2, P_1_1);
	wire S_3_0_3;
	wire C_3_0_3;
	fullAdder FA_3_0_3(S_3_0_3, C_3_0_3, S_2_0_3,  P_2_1, P_3_0);
	wire S_3_0_4;
	wire C_3_0_4;
	fullAdder FA_3_0_4(S_3_0_4, C_3_0_4, C_2_0_3,  S_2_0_4, P_4_0);
	wire S_3_0_5;
	wire C_3_0_5;
	fullAdder FA_3_0_5(S_3_0_5, C_3_0_5, C_2_0_4,  S_2_0_5, P_5_0);
	wire S_3_0_6;
	wire C_3_0_6;
	fullAdder FA_3_0_6(S_3_0_6, C_3_0_6, C_2_0_5,  S_2_0_6, S_1_3_6);
	wire S_3_0_7;
	wire C_3_0_7;
	fullAdder FA_3_0_7(S_3_0_7, C_3_0_7, C_2_0_6,  S_2_0_7, S_1_3_7);
	wire S_3_0_8;
	wire C_3_0_8;
	fullAdder FA_3_0_8(S_3_0_8, C_3_0_8, C_2_0_7,  S_2_0_8, S_1_3_8);
	wire S_3_0_9;
	wire C_3_0_9;
	fullAdder FA_3_0_9(S_3_0_9, C_3_0_9, C_2_0_8,  S_2_0_9, S_1_3_9);
	wire S_3_0_10;
	wire C_3_0_10;
	fullAdder FA_3_0_10(S_3_0_10, C_3_0_10, C_2_0_9,  S_2_0_10, S_1_3_10);
	wire S_3_0_11;
	wire C_3_0_11;
	fullAdder FA_3_0_11(S_3_0_11, C_3_0_11, C_2_0_10,  S_2_0_11, P_7_4);
	wire S_3_0_12;
	wire C_3_0_12;
	fullAdder FA_3_0_12(S_3_0_12, C_3_0_12, C_2_0_11,  S_2_0_12, C_1_0_11);
	wire S_3_0_13;
	wire C_3_0_13;
	fullAdder FA_3_0_13(S_3_0_13, C_3_0_13, P_6_7,  P_7_6, C_2_0_12);

	wire [13:0] in1 = {P_7_7, S_3_0_13, S_3_0_12, S_3_0_11, S_3_0_10, S_3_0_9, S_3_0_8, S_3_0_7, S_3_0_6, S_3_0_5, S_3_0_4, S_3_0_3, S_3_0_2, P_0_1};
	wire [13:0] in2 = {C_3_0_13, C_3_0_12, C_3_0_11, C_3_0_10, C_3_0_9, C_3_0_8, C_3_0_7, C_3_0_6, C_3_0_5, C_3_0_4, C_3_0_3, C_3_0_2, P_2_0, P_1_0};

	wire [14:0] ans;
	assign ans = in1 + in2;
	assign out = {ans, P_0_0};

	endmodule;
module wallace8_orig(out, a, b);

	input [15:0] a;
	input [15:0] b;
	output [31:0] out;


	wire P_0_0;
	wire P_0_1;
	wire P_0_2;
	wire P_0_3;
	wire P_0_4;
	wire P_0_5;
	wire P_0_6;
	wire P_0_7;
	wire P_0_8;
	wire P_0_9;
	wire P_0_10;
	wire P_0_11;
	wire P_0_12;
	wire P_0_13;
	wire P_0_14;
	wire P_0_15;
	wire P_1_0;
	wire P_1_1;
	wire P_1_2;
	wire P_1_3;
	wire P_1_4;
	wire P_1_5;
	wire P_1_6;
	wire P_1_7;
	wire P_1_8;
	wire P_1_9;
	wire P_1_10;
	wire P_1_11;
	wire P_1_12;
	wire P_1_13;
	wire P_1_14;
	wire P_1_15;
	wire P_2_0;
	wire P_2_1;
	wire P_2_2;
	wire P_2_3;
	wire P_2_4;
	wire P_2_5;
	wire P_2_6;
	wire P_2_7;
	wire P_2_8;
	wire P_2_9;
	wire P_2_10;
	wire P_2_11;
	wire P_2_12;
	wire P_2_13;
	wire P_2_14;
	wire P_2_15;
	wire P_3_0;
	wire P_3_1;
	wire P_3_2;
	wire P_3_3;
	wire P_3_4;
	wire P_3_5;
	wire P_3_6;
	wire P_3_7;
	wire P_3_8;
	wire P_3_9;
	wire P_3_10;
	wire P_3_11;
	wire P_3_12;
	wire P_3_13;
	wire P_3_14;
	wire P_3_15;
	wire P_4_0;
	wire P_4_1;
	wire P_4_2;
	wire P_4_3;
	wire P_4_4;
	wire P_4_5;
	wire P_4_6;
	wire P_4_7;
	wire P_4_8;
	wire P_4_9;
	wire P_4_10;
	wire P_4_11;
	wire P_4_12;
	wire P_4_13;
	wire P_4_14;
	wire P_4_15;
	wire P_5_0;
	wire P_5_1;
	wire P_5_2;
	wire P_5_3;
	wire P_5_4;
	wire P_5_5;
	wire P_5_6;
	wire P_5_7;
	wire P_5_8;
	wire P_5_9;
	wire P_5_10;
	wire P_5_11;
	wire P_5_12;
	wire P_5_13;
	wire P_5_14;
	wire P_5_15;
	wire P_6_0;
	wire P_6_1;
	wire P_6_2;
	wire P_6_3;
	wire P_6_4;
	wire P_6_5;
	wire P_6_6;
	wire P_6_7;
	wire P_6_8;
	wire P_6_9;
	wire P_6_10;
	wire P_6_11;
	wire P_6_12;
	wire P_6_13;
	wire P_6_14;
	wire P_6_15;
	wire P_7_0;
	wire P_7_1;
	wire P_7_2;
	wire P_7_3;
	wire P_7_4;
	wire P_7_5;
	wire P_7_6;
	wire P_7_7;
	wire P_7_8;
	wire P_7_9;
	wire P_7_10;
	wire P_7_11;
	wire P_7_12;
	wire P_7_13;
	wire P_7_14;
	wire P_7_15;
	wire P_8_0;
	wire P_8_1;
	wire P_8_2;
	wire P_8_3;
	wire P_8_4;
	wire P_8_5;
	wire P_8_6;
	wire P_8_7;
	wire P_8_8;
	wire P_8_9;
	wire P_8_10;
	wire P_8_11;
	wire P_8_12;
	wire P_8_13;
	wire P_8_14;
	wire P_8_15;
	wire P_9_0;
	wire P_9_1;
	wire P_9_2;
	wire P_9_3;
	wire P_9_4;
	wire P_9_5;
	wire P_9_6;
	wire P_9_7;
	wire P_9_8;
	wire P_9_9;
	wire P_9_10;
	wire P_9_11;
	wire P_9_12;
	wire P_9_13;
	wire P_9_14;
	wire P_9_15;
	wire P_10_0;
	wire P_10_1;
	wire P_10_2;
	wire P_10_3;
	wire P_10_4;
	wire P_10_5;
	wire P_10_6;
	wire P_10_7;
	wire P_10_8;
	wire P_10_9;
	wire P_10_10;
	wire P_10_11;
	wire P_10_12;
	wire P_10_13;
	wire P_10_14;
	wire P_10_15;
	wire P_11_0;
	wire P_11_1;
	wire P_11_2;
	wire P_11_3;
	wire P_11_4;
	wire P_11_5;
	wire P_11_6;
	wire P_11_7;
	wire P_11_8;
	wire P_11_9;
	wire P_11_10;
	wire P_11_11;
	wire P_11_12;
	wire P_11_13;
	wire P_11_14;
	wire P_11_15;
	wire P_12_0;
	wire P_12_1;
	wire P_12_2;
	wire P_12_3;
	wire P_12_4;
	wire P_12_5;
	wire P_12_6;
	wire P_12_7;
	wire P_12_8;
	wire P_12_9;
	wire P_12_10;
	wire P_12_11;
	wire P_12_12;
	wire P_12_13;
	wire P_12_14;
	wire P_12_15;
	wire P_13_0;
	wire P_13_1;
	wire P_13_2;
	wire P_13_3;
	wire P_13_4;
	wire P_13_5;
	wire P_13_6;
	wire P_13_7;
	wire P_13_8;
	wire P_13_9;
	wire P_13_10;
	wire P_13_11;
	wire P_13_12;
	wire P_13_13;
	wire P_13_14;
	wire P_13_15;
	wire P_14_0;
	wire P_14_1;
	wire P_14_2;
	wire P_14_3;
	wire P_14_4;
	wire P_14_5;
	wire P_14_6;
	wire P_14_7;
	wire P_14_8;
	wire P_14_9;
	wire P_14_10;
	wire P_14_11;
	wire P_14_12;
	wire P_14_13;
	wire P_14_14;
	wire P_14_15;
	wire P_15_0;
	wire P_15_1;
	wire P_15_2;
	wire P_15_3;
	wire P_15_4;
	wire P_15_5;
	wire P_15_6;
	wire P_15_7;
	wire P_15_8;
	wire P_15_9;
	wire P_15_10;
	wire P_15_11;
	wire P_15_12;
	wire P_15_13;
	wire P_15_14;
	wire P_15_15;
 /************************** AND gate DOT PRODUCT matrix ********************************/ 
	and A00(P_0_0, a[0], b[0]);
	and A01(P_0_1, a[0], b[1]);
	and A02(P_0_2, a[0], b[2]);
	and A03(P_0_3, a[0], b[3]);
	and A04(P_0_4, a[0], b[4]);
	and A05(P_0_5, a[0], b[5]);
	and A06(P_0_6, a[0], b[6]);
	and A07(P_0_7, a[0], b[7]);
	and A08(P_0_8, a[0], b[8]);
	and A09(P_0_9, a[0], b[9]);
	and A010(P_0_10, a[0], b[10]);
	and A011(P_0_11, a[0], b[11]);
	and A012(P_0_12, a[0], b[12]);
	and A013(P_0_13, a[0], b[13]);
	and A014(P_0_14, a[0], b[14]);
	and A015(P_0_15, a[0], b[15]);
	and A10(P_1_0, a[1], b[0]);
	and A11(P_1_1, a[1], b[1]);
	and A12(P_1_2, a[1], b[2]);
	and A13(P_1_3, a[1], b[3]);
	and A14(P_1_4, a[1], b[4]);
	and A15(P_1_5, a[1], b[5]);
	and A16(P_1_6, a[1], b[6]);
	and A17(P_1_7, a[1], b[7]);
	and A18(P_1_8, a[1], b[8]);
	and A19(P_1_9, a[1], b[9]);
	and A110(P_1_10, a[1], b[10]);
	and A111(P_1_11, a[1], b[11]);
	and A112(P_1_12, a[1], b[12]);
	and A113(P_1_13, a[1], b[13]);
	and A114(P_1_14, a[1], b[14]);
	and A115(P_1_15, a[1], b[15]);
	and A20(P_2_0, a[2], b[0]);
	and A21(P_2_1, a[2], b[1]);
	and A22(P_2_2, a[2], b[2]);
	and A23(P_2_3, a[2], b[3]);
	and A24(P_2_4, a[2], b[4]);
	and A25(P_2_5, a[2], b[5]);
	and A26(P_2_6, a[2], b[6]);
	and A27(P_2_7, a[2], b[7]);
	and A28(P_2_8, a[2], b[8]);
	and A29(P_2_9, a[2], b[9]);
	and A210(P_2_10, a[2], b[10]);
	and A211(P_2_11, a[2], b[11]);
	and A212(P_2_12, a[2], b[12]);
	and A213(P_2_13, a[2], b[13]);
	and A214(P_2_14, a[2], b[14]);
	and A215(P_2_15, a[2], b[15]);
	and A30(P_3_0, a[3], b[0]);
	and A31(P_3_1, a[3], b[1]);
	and A32(P_3_2, a[3], b[2]);
	and A33(P_3_3, a[3], b[3]);
	and A34(P_3_4, a[3], b[4]);
	and A35(P_3_5, a[3], b[5]);
	and A36(P_3_6, a[3], b[6]);
	and A37(P_3_7, a[3], b[7]);
	and A38(P_3_8, a[3], b[8]);
	and A39(P_3_9, a[3], b[9]);
	and A310(P_3_10, a[3], b[10]);
	and A311(P_3_11, a[3], b[11]);
	and A312(P_3_12, a[3], b[12]);
	and A313(P_3_13, a[3], b[13]);
	and A314(P_3_14, a[3], b[14]);
	and A315(P_3_15, a[3], b[15]);
	and A40(P_4_0, a[4], b[0]);
	and A41(P_4_1, a[4], b[1]);
	and A42(P_4_2, a[4], b[2]);
	and A43(P_4_3, a[4], b[3]);
	and A44(P_4_4, a[4], b[4]);
	and A45(P_4_5, a[4], b[5]);
	and A46(P_4_6, a[4], b[6]);
	and A47(P_4_7, a[4], b[7]);
	and A48(P_4_8, a[4], b[8]);
	and A49(P_4_9, a[4], b[9]);
	and A410(P_4_10, a[4], b[10]);
	and A411(P_4_11, a[4], b[11]);
	and A412(P_4_12, a[4], b[12]);
	and A413(P_4_13, a[4], b[13]);
	and A414(P_4_14, a[4], b[14]);
	and A415(P_4_15, a[4], b[15]);
	and A50(P_5_0, a[5], b[0]);
	and A51(P_5_1, a[5], b[1]);
	and A52(P_5_2, a[5], b[2]);
	and A53(P_5_3, a[5], b[3]);
	and A54(P_5_4, a[5], b[4]);
	and A55(P_5_5, a[5], b[5]);
	and A56(P_5_6, a[5], b[6]);
	and A57(P_5_7, a[5], b[7]);
	and A58(P_5_8, a[5], b[8]);
	and A59(P_5_9, a[5], b[9]);
	and A510(P_5_10, a[5], b[10]);
	and A511(P_5_11, a[5], b[11]);
	and A512(P_5_12, a[5], b[12]);
	and A513(P_5_13, a[5], b[13]);
	and A514(P_5_14, a[5], b[14]);
	and A515(P_5_15, a[5], b[15]);
	and A60(P_6_0, a[6], b[0]);
	and A61(P_6_1, a[6], b[1]);
	and A62(P_6_2, a[6], b[2]);
	and A63(P_6_3, a[6], b[3]);
	and A64(P_6_4, a[6], b[4]);
	and A65(P_6_5, a[6], b[5]);
	and A66(P_6_6, a[6], b[6]);
	and A67(P_6_7, a[6], b[7]);
	and A68(P_6_8, a[6], b[8]);
	and A69(P_6_9, a[6], b[9]);
	and A610(P_6_10, a[6], b[10]);
	and A611(P_6_11, a[6], b[11]);
	and A612(P_6_12, a[6], b[12]);
	and A613(P_6_13, a[6], b[13]);
	and A614(P_6_14, a[6], b[14]);
	and A615(P_6_15, a[6], b[15]);
	and A70(P_7_0, a[7], b[0]);
	and A71(P_7_1, a[7], b[1]);
	and A72(P_7_2, a[7], b[2]);
	and A73(P_7_3, a[7], b[3]);
	and A74(P_7_4, a[7], b[4]);
	and A75(P_7_5, a[7], b[5]);
	and A76(P_7_6, a[7], b[6]);
	and A77(P_7_7, a[7], b[7]);
	and A78(P_7_8, a[7], b[8]);
	and A79(P_7_9, a[7], b[9]);
	and A710(P_7_10, a[7], b[10]);
	and A711(P_7_11, a[7], b[11]);
	and A712(P_7_12, a[7], b[12]);
	and A713(P_7_13, a[7], b[13]);
	and A714(P_7_14, a[7], b[14]);
	and A715(P_7_15, a[7], b[15]);
	and A80(P_8_0, a[8], b[0]);
	and A81(P_8_1, a[8], b[1]);
	and A82(P_8_2, a[8], b[2]);
	and A83(P_8_3, a[8], b[3]);
	and A84(P_8_4, a[8], b[4]);
	and A85(P_8_5, a[8], b[5]);
	and A86(P_8_6, a[8], b[6]);
	and A87(P_8_7, a[8], b[7]);
	and A88(P_8_8, a[8], b[8]);
	and A89(P_8_9, a[8], b[9]);
	and A810(P_8_10, a[8], b[10]);
	and A811(P_8_11, a[8], b[11]);
	and A812(P_8_12, a[8], b[12]);
	and A813(P_8_13, a[8], b[13]);
	and A814(P_8_14, a[8], b[14]);
	and A815(P_8_15, a[8], b[15]);
	and A90(P_9_0, a[9], b[0]);
	and A91(P_9_1, a[9], b[1]);
	and A92(P_9_2, a[9], b[2]);
	and A93(P_9_3, a[9], b[3]);
	and A94(P_9_4, a[9], b[4]);
	and A95(P_9_5, a[9], b[5]);
	and A96(P_9_6, a[9], b[6]);
	and A97(P_9_7, a[9], b[7]);
	and A98(P_9_8, a[9], b[8]);
	and A99(P_9_9, a[9], b[9]);
	and A910(P_9_10, a[9], b[10]);
	and A911(P_9_11, a[9], b[11]);
	and A912(P_9_12, a[9], b[12]);
	and A913(P_9_13, a[9], b[13]);
	and A914(P_9_14, a[9], b[14]);
	and A915(P_9_15, a[9], b[15]);
	and A100(P_10_0, a[10], b[0]);
	and A101(P_10_1, a[10], b[1]);
	and A102(P_10_2, a[10], b[2]);
	and A103(P_10_3, a[10], b[3]);
	and A104(P_10_4, a[10], b[4]);
	and A105(P_10_5, a[10], b[5]);
	and A106(P_10_6, a[10], b[6]);
	and A107(P_10_7, a[10], b[7]);
	and A108(P_10_8, a[10], b[8]);
	and A109(P_10_9, a[10], b[9]);
	and A1010(P_10_10, a[10], b[10]);
	and A1011(P_10_11, a[10], b[11]);
	and A1012(P_10_12, a[10], b[12]);
	and A1013(P_10_13, a[10], b[13]);
	and A1014(P_10_14, a[10], b[14]);
	and A1015(P_10_15, a[10], b[15]);
	and A110(P_11_0, a[11], b[0]);
	and A111(P_11_1, a[11], b[1]);
	and A112(P_11_2, a[11], b[2]);
	and A113(P_11_3, a[11], b[3]);
	and A114(P_11_4, a[11], b[4]);
	and A115(P_11_5, a[11], b[5]);
	and A116(P_11_6, a[11], b[6]);
	and A117(P_11_7, a[11], b[7]);
	and A118(P_11_8, a[11], b[8]);
	and A119(P_11_9, a[11], b[9]);
	and A1110(P_11_10, a[11], b[10]);
	and A1111(P_11_11, a[11], b[11]);
	and A1112(P_11_12, a[11], b[12]);
	and A1113(P_11_13, a[11], b[13]);
	and A1114(P_11_14, a[11], b[14]);
	and A1115(P_11_15, a[11], b[15]);
	and A120(P_12_0, a[12], b[0]);
	and A121(P_12_1, a[12], b[1]);
	and A122(P_12_2, a[12], b[2]);
	and A123(P_12_3, a[12], b[3]);
	and A124(P_12_4, a[12], b[4]);
	and A125(P_12_5, a[12], b[5]);
	and A126(P_12_6, a[12], b[6]);
	and A127(P_12_7, a[12], b[7]);
	and A128(P_12_8, a[12], b[8]);
	and A129(P_12_9, a[12], b[9]);
	and A1210(P_12_10, a[12], b[10]);
	and A1211(P_12_11, a[12], b[11]);
	and A1212(P_12_12, a[12], b[12]);
	and A1213(P_12_13, a[12], b[13]);
	and A1214(P_12_14, a[12], b[14]);
	and A1215(P_12_15, a[12], b[15]);
	and A130(P_13_0, a[13], b[0]);
	and A131(P_13_1, a[13], b[1]);
	and A132(P_13_2, a[13], b[2]);
	and A133(P_13_3, a[13], b[3]);
	and A134(P_13_4, a[13], b[4]);
	and A135(P_13_5, a[13], b[5]);
	and A136(P_13_6, a[13], b[6]);
	and A137(P_13_7, a[13], b[7]);
	and A138(P_13_8, a[13], b[8]);
	and A139(P_13_9, a[13], b[9]);
	and A1310(P_13_10, a[13], b[10]);
	and A1311(P_13_11, a[13], b[11]);
	and A1312(P_13_12, a[13], b[12]);
	and A1313(P_13_13, a[13], b[13]);
	and A1314(P_13_14, a[13], b[14]);
	and A1315(P_13_15, a[13], b[15]);
	and A140(P_14_0, a[14], b[0]);
	and A141(P_14_1, a[14], b[1]);
	and A142(P_14_2, a[14], b[2]);
	and A143(P_14_3, a[14], b[3]);
	and A144(P_14_4, a[14], b[4]);
	and A145(P_14_5, a[14], b[5]);
	and A146(P_14_6, a[14], b[6]);
	and A147(P_14_7, a[14], b[7]);
	and A148(P_14_8, a[14], b[8]);
	and A149(P_14_9, a[14], b[9]);
	and A1410(P_14_10, a[14], b[10]);
	and A1411(P_14_11, a[14], b[11]);
	and A1412(P_14_12, a[14], b[12]);
	and A1413(P_14_13, a[14], b[13]);
	and A1414(P_14_14, a[14], b[14]);
	and A1415(P_14_15, a[14], b[15]);
	and A150(P_15_0, a[15], b[0]);
	and A151(P_15_1, a[15], b[1]);
	and A152(P_15_2, a[15], b[2]);
	and A153(P_15_3, a[15], b[3]);
	and A154(P_15_4, a[15], b[4]);
	and A155(P_15_5, a[15], b[5]);
	and A156(P_15_6, a[15], b[6]);
	and A157(P_15_7, a[15], b[7]);
	and A158(P_15_8, a[15], b[8]);
	and A159(P_15_9, a[15], b[9]);
	and A1510(P_15_10, a[15], b[10]);
	and A1511(P_15_11, a[15], b[11]);
	and A1512(P_15_12, a[15], b[12]);
	and A1513(P_15_13, a[15], b[13]);
	and A1514(P_15_14, a[15], b[14]);
	and A1515(P_15_15, a[15], b[15]);
	wire S_0_1_0_1;
	wire C_0_1_0_1;
	wire S_0_1_0_2;
	wire C_0_1_0_2;
	wire S_0_1_0_3;
	wire C_0_1_0_3;
	wire S_0_1_0_4;
	wire C_0_1_0_4;
	wire S_0_1_0_5;
	wire C_0_1_0_5;
	wire S_0_1_0_6;
	wire C_0_1_0_6;
	wire S_0_1_0_7;
	wire C_0_1_0_7;
	wire S_0_1_0_8;
	wire C_0_1_0_8;
	wire S_0_1_0_9;
	wire C_0_1_0_9;
	wire S_0_1_0_10;
	wire C_0_1_0_10;
	wire S_0_1_0_11;
	wire C_0_1_0_11;
	wire S_0_1_0_12;
	wire C_0_1_0_12;
	wire S_0_1_0_13;
	wire C_0_1_0_13;
	wire S_0_1_0_14;
	wire C_0_1_0_14;
	wire S_0_1_0_15;
	wire C_0_1_0_15;
	wire S_0_1_0_16;
	wire C_0_1_0_16;
	wire S_0_2_3_4;
	wire C_0_2_3_4;
	wire S_0_2_3_5;
	wire C_0_2_3_5;
	wire S_0_2_3_6;
	wire C_0_2_3_6;
	wire S_0_2_3_7;
	wire C_0_2_3_7;
	wire S_0_2_3_8;
	wire C_0_2_3_8;
	wire S_0_2_3_9;
	wire C_0_2_3_9;
	wire S_0_2_3_10;
	wire C_0_2_3_10;
	wire S_0_2_3_11;
	wire C_0_2_3_11;
	wire S_0_2_3_12;
	wire C_0_2_3_12;
	wire S_0_2_3_13;
	wire C_0_2_3_13;
	wire S_0_2_3_14;
	wire C_0_2_3_14;
	wire S_0_2_3_15;
	wire C_0_2_3_15;
	wire S_0_2_3_16;
	wire C_0_2_3_16;
	wire S_0_2_3_17;
	wire C_0_2_3_17;
	wire S_0_2_3_18;
	wire C_0_2_3_18;
	wire S_0_2_3_19;
	wire C_0_2_3_19;
	wire S_0_3_6_7;
	wire C_0_3_6_7;
	wire S_0_3_6_8;
	wire C_0_3_6_8;
	wire S_0_3_6_9;
	wire C_0_3_6_9;
	wire S_0_3_6_10;
	wire C_0_3_6_10;
	wire S_0_3_6_11;
	wire C_0_3_6_11;
	wire S_0_3_6_12;
	wire C_0_3_6_12;
	wire S_0_3_6_13;
	wire C_0_3_6_13;
	wire S_0_3_6_14;
	wire C_0_3_6_14;
	wire S_0_3_6_15;
	wire C_0_3_6_15;
	wire S_0_3_6_16;
	wire C_0_3_6_16;
	wire S_0_3_6_17;
	wire C_0_3_6_17;
	wire S_0_3_6_18;
	wire C_0_3_6_18;
	wire S_0_3_6_19;
	wire C_0_3_6_19;
	wire S_0_3_6_20;
	wire C_0_3_6_20;
	wire S_0_3_6_21;
	wire C_0_3_6_21;
	wire S_0_3_6_22;
	wire C_0_3_6_22;
	wire S_0_4_9_10;
	wire C_0_4_9_10;
	wire S_0_4_9_11;
	wire C_0_4_9_11;
	wire S_0_4_9_12;
	wire C_0_4_9_12;
	wire S_0_4_9_13;
	wire C_0_4_9_13;
	wire S_0_4_9_14;
	wire C_0_4_9_14;
	wire S_0_4_9_15;
	wire C_0_4_9_15;
	wire S_0_4_9_16;
	wire C_0_4_9_16;
	wire S_0_4_9_17;
	wire C_0_4_9_17;
	wire S_0_4_9_18;
	wire C_0_4_9_18;
	wire S_0_4_9_19;
	wire C_0_4_9_19;
	wire S_0_4_9_20;
	wire C_0_4_9_20;
	wire S_0_4_9_21;
	wire C_0_4_9_21;
	wire S_0_4_9_22;
	wire C_0_4_9_22;
	wire S_0_4_9_23;
	wire C_0_4_9_23;
	wire S_0_4_9_24;
	wire C_0_4_9_24;
	wire S_0_4_9_25;
	wire C_0_4_9_25;
	wire S_0_5_12_13;
	wire C_0_5_12_13;
	wire S_0_5_12_14;
	wire C_0_5_12_14;
	wire S_0_5_12_15;
	wire C_0_5_12_15;
	wire S_0_5_12_16;
	wire C_0_5_12_16;
	wire S_0_5_12_17;
	wire C_0_5_12_17;
	wire S_0_5_12_18;
	wire C_0_5_12_18;
	wire S_0_5_12_19;
	wire C_0_5_12_19;
	wire S_0_5_12_20;
	wire C_0_5_12_20;
	wire S_0_5_12_21;
	wire C_0_5_12_21;
	wire S_0_5_12_22;
	wire C_0_5_12_22;
	wire S_0_5_12_23;
	wire C_0_5_12_23;
	wire S_0_5_12_24;
	wire C_0_5_12_24;
	wire S_0_5_12_25;
	wire C_0_5_12_25;
	wire S_0_5_12_26;
	wire C_0_5_12_26;
	wire S_0_5_12_27;
	wire C_0_5_12_27;
	wire S_0_5_12_28;
	wire C_0_5_12_28;
	wire S_1_1_0_2;
	wire C_1_1_0_2;
	wire S_1_1_0_3;
	wire C_1_1_0_3;
	wire S_1_1_0_4;
	wire C_1_1_0_4;
	wire S_1_1_0_5;
	wire C_1_1_0_5;
	wire S_1_1_0_6;
	wire C_1_1_0_6;
	wire S_1_1_0_7;
	wire C_1_1_0_7;
	wire S_1_1_0_8;
	wire C_1_1_0_8;
	wire S_1_1_0_9;
	wire C_1_1_0_9;
	wire S_1_1_0_10;
	wire C_1_1_0_10;
	wire S_1_1_0_11;
	wire C_1_1_0_11;
	wire S_1_1_0_12;
	wire C_1_1_0_12;
	wire S_1_1_0_13;
	wire C_1_1_0_13;
	wire S_1_1_0_14;
	wire C_1_1_0_14;
	wire S_1_1_0_15;
	wire C_1_1_0_15;
	wire S_1_1_0_16;
	wire C_1_1_0_16;
	wire S_1_1_0_17;
	wire C_1_1_0_17;
	wire S_1_2_3_6;
	wire C_1_2_3_6;
	wire S_1_2_3_7;
	wire C_1_2_3_7;
	wire S_1_2_3_8;
	wire C_1_2_3_8;
	wire S_1_2_3_9;
	wire C_1_2_3_9;
	wire S_1_2_3_10;
	wire C_1_2_3_10;
	wire S_1_2_3_11;
	wire C_1_2_3_11;
	wire S_1_2_3_12;
	wire C_1_2_3_12;
	wire S_1_2_3_13;
	wire C_1_2_3_13;
	wire S_1_2_3_14;
	wire C_1_2_3_14;
	wire S_1_2_3_15;
	wire C_1_2_3_15;
	wire S_1_2_3_16;
	wire C_1_2_3_16;
	wire S_1_2_3_17;
	wire C_1_2_3_17;
	wire S_1_2_3_18;
	wire C_1_2_3_18;
	wire S_1_2_3_19;
	wire C_1_2_3_19;
	wire S_1_2_3_20;
	wire C_1_2_3_20;
	wire S_1_2_3_21;
	wire C_1_2_3_21;
	wire S_1_2_3_22;
	wire C_1_2_3_22;
	wire S_1_2_3_23;
	wire C_1_2_3_23;
	wire S_1_3_6_11;
	wire C_1_3_6_11;
	wire S_1_3_6_12;
	wire C_1_3_6_12;
	wire S_1_3_6_13;
	wire C_1_3_6_13;
	wire S_1_3_6_14;
	wire C_1_3_6_14;
	wire S_1_3_6_15;
	wire C_1_3_6_15;
	wire S_1_3_6_16;
	wire C_1_3_6_16;
	wire S_1_3_6_17;
	wire C_1_3_6_17;
	wire S_1_3_6_18;
	wire C_1_3_6_18;
	wire S_1_3_6_19;
	wire C_1_3_6_19;
	wire S_1_3_6_20;
	wire C_1_3_6_20;
	wire S_1_3_6_21;
	wire C_1_3_6_21;
	wire S_1_3_6_22;
	wire C_1_3_6_22;
	wire S_1_3_6_23;
	wire C_1_3_6_23;
	wire S_1_3_6_24;
	wire C_1_3_6_24;
	wire S_1_3_6_25;
	wire C_1_3_6_25;
	wire S_1_3_6_26;
	wire C_1_3_6_26;
	wire S_2_1_0_3;
	wire C_2_1_0_3;
	wire S_2_1_0_4;
	wire C_2_1_0_4;
	wire S_2_1_0_5;
	wire C_2_1_0_5;
	wire S_2_1_0_6;
	wire C_2_1_0_6;
	wire S_2_1_0_7;
	wire C_2_1_0_7;
	wire S_2_1_0_8;
	wire C_2_1_0_8;
	wire S_2_1_0_9;
	wire C_2_1_0_9;
	wire S_2_1_0_10;
	wire C_2_1_0_10;
	wire S_2_1_0_11;
	wire C_2_1_0_11;
	wire S_2_1_0_12;
	wire C_2_1_0_12;
	wire S_2_1_0_13;
	wire C_2_1_0_13;
	wire S_2_1_0_14;
	wire C_2_1_0_14;
	wire S_2_1_0_15;
	wire C_2_1_0_15;
	wire S_2_1_0_16;
	wire C_2_1_0_16;
	wire S_2_1_0_17;
	wire C_2_1_0_17;
	wire S_2_1_0_18;
	wire C_2_1_0_18;
	wire S_2_1_0_19;
	wire C_2_1_0_19;
	wire S_2_1_0_20;
	wire C_2_1_0_20;
	wire S_2_2_3_9;
	wire C_2_2_3_9;
	wire S_2_2_3_10;
	wire C_2_2_3_10;
	wire S_2_2_3_11;
	wire C_2_2_3_11;
	wire S_2_2_3_12;
	wire C_2_2_3_12;
	wire S_2_2_3_13;
	wire C_2_2_3_13;
	wire S_2_2_3_14;
	wire C_2_2_3_14;
	wire S_2_2_3_15;
	wire C_2_2_3_15;
	wire S_2_2_3_16;
	wire C_2_2_3_16;
	wire S_2_2_3_17;
	wire C_2_2_3_17;
	wire S_2_2_3_18;
	wire C_2_2_3_18;
	wire S_2_2_3_19;
	wire C_2_2_3_19;
	wire S_2_2_3_20;
	wire C_2_2_3_20;
	wire S_2_2_3_21;
	wire C_2_2_3_21;
	wire S_2_2_3_22;
	wire C_2_2_3_22;
	wire S_2_2_3_23;
	wire C_2_2_3_23;
	wire S_2_2_3_24;
	wire C_2_2_3_24;
	wire S_2_2_3_25;
	wire C_2_2_3_25;
	wire S_2_2_3_26;
	wire C_2_2_3_26;
	wire S_2_2_3_27;
	wire C_2_2_3_27;
	wire S_3_1_0_4;
	wire C_3_1_0_4;
	wire S_3_1_0_5;
	wire C_3_1_0_5;
	wire S_3_1_0_6;
	wire C_3_1_0_6;
	wire S_3_1_0_7;
	wire C_3_1_0_7;
	wire S_3_1_0_8;
	wire C_3_1_0_8;
	wire S_3_1_0_9;
	wire C_3_1_0_9;
	wire S_3_1_0_10;
	wire C_3_1_0_10;
	wire S_3_1_0_11;
	wire C_3_1_0_11;
	wire S_3_1_0_12;
	wire C_3_1_0_12;
	wire S_3_1_0_13;
	wire C_3_1_0_13;
	wire S_3_1_0_14;
	wire C_3_1_0_14;
	wire S_3_1_0_15;
	wire C_3_1_0_15;
	wire S_3_1_0_16;
	wire C_3_1_0_16;
	wire S_3_1_0_17;
	wire C_3_1_0_17;
	wire S_3_1_0_18;
	wire C_3_1_0_18;
	wire S_3_1_0_19;
	wire C_3_1_0_19;
	wire S_3_1_0_20;
	wire C_3_1_0_20;
	wire S_3_1_0_21;
	wire C_3_1_0_21;
	wire S_3_1_0_22;
	wire C_3_1_0_22;
	wire S_3_1_0_23;
	wire C_3_1_0_23;
	wire S_4_1_0_5;
	wire C_4_1_0_5;
	wire S_4_1_0_6;
	wire C_4_1_0_6;
	wire S_4_1_0_7;
	wire C_4_1_0_7;
	wire S_4_1_0_8;
	wire C_4_1_0_8;
	wire S_4_1_0_9;
	wire C_4_1_0_9;
	wire S_4_1_0_10;
	wire C_4_1_0_10;
	wire S_4_1_0_11;
	wire C_4_1_0_11;
	wire S_4_1_0_12;
	wire C_4_1_0_12;
	wire S_4_1_0_13;
	wire C_4_1_0_13;
	wire S_4_1_0_14;
	wire C_4_1_0_14;
	wire S_4_1_0_15;
	wire C_4_1_0_15;
	wire S_4_1_0_16;
	wire C_4_1_0_16;
	wire S_4_1_0_17;
	wire C_4_1_0_17;
	wire S_4_1_0_18;
	wire C_4_1_0_18;
	wire S_4_1_0_19;
	wire C_4_1_0_19;
	wire S_4_1_0_20;
	wire C_4_1_0_20;
	wire S_4_1_0_21;
	wire C_4_1_0_21;
	wire S_4_1_0_22;
	wire C_4_1_0_22;
	wire S_4_1_0_23;
	wire C_4_1_0_23;
	wire S_4_1_0_24;
	wire C_4_1_0_24;
	wire S_4_1_0_25;
	wire C_4_1_0_25;
	wire S_4_1_0_26;
	wire C_4_1_0_26;
	wire S_4_1_0_27;
	wire C_4_1_0_27;
	wire S_4_1_0_28;
	wire C_4_1_0_28;
	wire S_5_1_0_6;
	wire C_5_1_0_6;
	wire S_5_1_0_7;
	wire C_5_1_0_7;
	wire S_5_1_0_8;
	wire C_5_1_0_8;
	wire S_5_1_0_9;
	wire C_5_1_0_9;
	wire S_5_1_0_10;
	wire C_5_1_0_10;
	wire S_5_1_0_11;
	wire C_5_1_0_11;
	wire S_5_1_0_12;
	wire C_5_1_0_12;
	wire S_5_1_0_13;
	wire C_5_1_0_13;
	wire S_5_1_0_14;
	wire C_5_1_0_14;
	wire S_5_1_0_15;
	wire C_5_1_0_15;
	wire S_5_1_0_16;
	wire C_5_1_0_16;
	wire S_5_1_0_17;
	wire C_5_1_0_17;
	wire S_5_1_0_18;
	wire C_5_1_0_18;
	wire S_5_1_0_19;
	wire C_5_1_0_19;
	wire S_5_1_0_20;
	wire C_5_1_0_20;
	wire S_5_1_0_21;
	wire C_5_1_0_21;
	wire S_5_1_0_22;
	wire C_5_1_0_22;
	wire S_5_1_0_23;
	wire C_5_1_0_23;
	wire S_5_1_0_24;
	wire C_5_1_0_24;
	wire S_5_1_0_25;
	wire C_5_1_0_25;
	wire S_5_1_0_26;
	wire C_5_1_0_26;
	wire S_5_1_0_27;
	wire C_5_1_0_27;
	wire S_5_1_0_28;
	wire C_5_1_0_28;
	wire S_5_1_0_29;
	wire C_5_1_0_29;
 /************************** Height - 0 ********************************/ 
 /************************** Layer - 0 ********************************/ 
	halfAdder HA_0_1_0_1(S_0_1_0_1, C_0_1_0_1, P_0_1, P_1_0);
	fullAdder FA_0_1_0_2(S_0_1_0_2, C_0_1_0_2, P_0_2, P_1_1, P_2_0);
	fullAdder FA_0_1_0_3(S_0_1_0_3, C_0_1_0_3, P_0_3, P_1_2, P_2_1);
	fullAdder FA_0_1_0_4(S_0_1_0_4, C_0_1_0_4, P_0_4, P_1_3, P_2_2);
	fullAdder FA_0_1_0_5(S_0_1_0_5, C_0_1_0_5, P_0_5, P_1_4, P_2_3);
	fullAdder FA_0_1_0_6(S_0_1_0_6, C_0_1_0_6, P_0_6, P_1_5, P_2_4);
	fullAdder FA_0_1_0_7(S_0_1_0_7, C_0_1_0_7, P_0_7, P_1_6, P_2_5);
	fullAdder FA_0_1_0_8(S_0_1_0_8, C_0_1_0_8, P_0_8, P_1_7, P_2_6);
	fullAdder FA_0_1_0_9(S_0_1_0_9, C_0_1_0_9, P_0_9, P_1_8, P_2_7);
	fullAdder FA_0_1_0_10(S_0_1_0_10, C_0_1_0_10, P_0_10, P_1_9, P_2_8);
	fullAdder FA_0_1_0_11(S_0_1_0_11, C_0_1_0_11, P_0_11, P_1_10, P_2_9);
	fullAdder FA_0_1_0_12(S_0_1_0_12, C_0_1_0_12, P_0_12, P_1_11, P_2_10);
	fullAdder FA_0_1_0_13(S_0_1_0_13, C_0_1_0_13, P_0_13, P_1_12, P_2_11);
	fullAdder FA_0_1_0_14(S_0_1_0_14, C_0_1_0_14, P_0_14, P_1_13, P_2_12);
	fullAdder FA_0_1_0_15(S_0_1_0_15, C_0_1_0_15, P_0_15, P_1_14, P_2_13);
	halfAdder HA_0_1_0_16(S_0_1_0_16, C_0_1_0_16, P_1_15, P_2_14);
 /************************** Layer - 3 ********************************/ 
	halfAdder HA_0_2_3_4(S_0_2_3_4, C_0_2_3_4, P_3_1, P_4_0);
	fullAdder FA_0_2_3_5(S_0_2_3_5, C_0_2_3_5, P_3_2, P_4_1, P_5_0);
	fullAdder FA_0_2_3_6(S_0_2_3_6, C_0_2_3_6, P_3_3, P_4_2, P_5_1);
	fullAdder FA_0_2_3_7(S_0_2_3_7, C_0_2_3_7, P_3_4, P_4_3, P_5_2);
	fullAdder FA_0_2_3_8(S_0_2_3_8, C_0_2_3_8, P_3_5, P_4_4, P_5_3);
	fullAdder FA_0_2_3_9(S_0_2_3_9, C_0_2_3_9, P_3_6, P_4_5, P_5_4);
	fullAdder FA_0_2_3_10(S_0_2_3_10, C_0_2_3_10, P_3_7, P_4_6, P_5_5);
	fullAdder FA_0_2_3_11(S_0_2_3_11, C_0_2_3_11, P_3_8, P_4_7, P_5_6);
	fullAdder FA_0_2_3_12(S_0_2_3_12, C_0_2_3_12, P_3_9, P_4_8, P_5_7);
	fullAdder FA_0_2_3_13(S_0_2_3_13, C_0_2_3_13, P_3_10, P_4_9, P_5_8);
	fullAdder FA_0_2_3_14(S_0_2_3_14, C_0_2_3_14, P_3_11, P_4_10, P_5_9);
	fullAdder FA_0_2_3_15(S_0_2_3_15, C_0_2_3_15, P_3_12, P_4_11, P_5_10);
	fullAdder FA_0_2_3_16(S_0_2_3_16, C_0_2_3_16, P_3_13, P_4_12, P_5_11);
	fullAdder FA_0_2_3_17(S_0_2_3_17, C_0_2_3_17, P_3_14, P_4_13, P_5_12);
	fullAdder FA_0_2_3_18(S_0_2_3_18, C_0_2_3_18, P_3_15, P_4_14, P_5_13);
	halfAdder HA_0_2_3_19(S_0_2_3_19, C_0_2_3_19, P_4_15, P_5_14);
 /************************** Layer - 6 ********************************/ 
	halfAdder HA_0_3_6_7(S_0_3_6_7, C_0_3_6_7, P_6_1, P_7_0);
	fullAdder FA_0_3_6_8(S_0_3_6_8, C_0_3_6_8, P_6_2, P_7_1, P_8_0);
	fullAdder FA_0_3_6_9(S_0_3_6_9, C_0_3_6_9, P_6_3, P_7_2, P_8_1);
	fullAdder FA_0_3_6_10(S_0_3_6_10, C_0_3_6_10, P_6_4, P_7_3, P_8_2);
	fullAdder FA_0_3_6_11(S_0_3_6_11, C_0_3_6_11, P_6_5, P_7_4, P_8_3);
	fullAdder FA_0_3_6_12(S_0_3_6_12, C_0_3_6_12, P_6_6, P_7_5, P_8_4);
	fullAdder FA_0_3_6_13(S_0_3_6_13, C_0_3_6_13, P_6_7, P_7_6, P_8_5);
	fullAdder FA_0_3_6_14(S_0_3_6_14, C_0_3_6_14, P_6_8, P_7_7, P_8_6);
	fullAdder FA_0_3_6_15(S_0_3_6_15, C_0_3_6_15, P_6_9, P_7_8, P_8_7);
	fullAdder FA_0_3_6_16(S_0_3_6_16, C_0_3_6_16, P_6_10, P_7_9, P_8_8);
	fullAdder FA_0_3_6_17(S_0_3_6_17, C_0_3_6_17, P_6_11, P_7_10, P_8_9);
	fullAdder FA_0_3_6_18(S_0_3_6_18, C_0_3_6_18, P_6_12, P_7_11, P_8_10);
	fullAdder FA_0_3_6_19(S_0_3_6_19, C_0_3_6_19, P_6_13, P_7_12, P_8_11);
	fullAdder FA_0_3_6_20(S_0_3_6_20, C_0_3_6_20, P_6_14, P_7_13, P_8_12);
	fullAdder FA_0_3_6_21(S_0_3_6_21, C_0_3_6_21, P_6_15, P_7_14, P_8_13);
	halfAdder HA_0_3_6_22(S_0_3_6_22, C_0_3_6_22, P_7_15, P_8_14);
 /************************** Layer - 9 ********************************/ 
	halfAdder HA_0_4_9_10(S_0_4_9_10, C_0_4_9_10, P_9_1, P_10_0);
	fullAdder FA_0_4_9_11(S_0_4_9_11, C_0_4_9_11, P_9_2, P_10_1, P_11_0);
	fullAdder FA_0_4_9_12(S_0_4_9_12, C_0_4_9_12, P_9_3, P_10_2, P_11_1);
	fullAdder FA_0_4_9_13(S_0_4_9_13, C_0_4_9_13, P_9_4, P_10_3, P_11_2);
	fullAdder FA_0_4_9_14(S_0_4_9_14, C_0_4_9_14, P_9_5, P_10_4, P_11_3);
	fullAdder FA_0_4_9_15(S_0_4_9_15, C_0_4_9_15, P_9_6, P_10_5, P_11_4);
	fullAdder FA_0_4_9_16(S_0_4_9_16, C_0_4_9_16, P_9_7, P_10_6, P_11_5);
	fullAdder FA_0_4_9_17(S_0_4_9_17, C_0_4_9_17, P_9_8, P_10_7, P_11_6);
	fullAdder FA_0_4_9_18(S_0_4_9_18, C_0_4_9_18, P_9_9, P_10_8, P_11_7);
	fullAdder FA_0_4_9_19(S_0_4_9_19, C_0_4_9_19, P_9_10, P_10_9, P_11_8);
	fullAdder FA_0_4_9_20(S_0_4_9_20, C_0_4_9_20, P_9_11, P_10_10, P_11_9);
	fullAdder FA_0_4_9_21(S_0_4_9_21, C_0_4_9_21, P_9_12, P_10_11, P_11_10);
	fullAdder FA_0_4_9_22(S_0_4_9_22, C_0_4_9_22, P_9_13, P_10_12, P_11_11);
	fullAdder FA_0_4_9_23(S_0_4_9_23, C_0_4_9_23, P_9_14, P_10_13, P_11_12);
	fullAdder FA_0_4_9_24(S_0_4_9_24, C_0_4_9_24, P_9_15, P_10_14, P_11_13);
	halfAdder HA_0_4_9_25(S_0_4_9_25, C_0_4_9_25, P_10_15, P_11_14);
 /************************** Layer - 12 ********************************/ 
	halfAdder HA_0_5_12_13(S_0_5_12_13, C_0_5_12_13, P_12_1, P_13_0);
	fullAdder FA_0_5_12_14(S_0_5_12_14, C_0_5_12_14, P_12_2, P_13_1, P_14_0);
	fullAdder FA_0_5_12_15(S_0_5_12_15, C_0_5_12_15, P_12_3, P_13_2, P_14_1);
	fullAdder FA_0_5_12_16(S_0_5_12_16, C_0_5_12_16, P_12_4, P_13_3, P_14_2);
	fullAdder FA_0_5_12_17(S_0_5_12_17, C_0_5_12_17, P_12_5, P_13_4, P_14_3);
	fullAdder FA_0_5_12_18(S_0_5_12_18, C_0_5_12_18, P_12_6, P_13_5, P_14_4);
	fullAdder FA_0_5_12_19(S_0_5_12_19, C_0_5_12_19, P_12_7, P_13_6, P_14_5);
	fullAdder FA_0_5_12_20(S_0_5_12_20, C_0_5_12_20, P_12_8, P_13_7, P_14_6);
	fullAdder FA_0_5_12_21(S_0_5_12_21, C_0_5_12_21, P_12_9, P_13_8, P_14_7);
	fullAdder FA_0_5_12_22(S_0_5_12_22, C_0_5_12_22, P_12_10, P_13_9, P_14_8);
	fullAdder FA_0_5_12_23(S_0_5_12_23, C_0_5_12_23, P_12_11, P_13_10, P_14_9);
	fullAdder FA_0_5_12_24(S_0_5_12_24, C_0_5_12_24, P_12_12, P_13_11, P_14_10);
	fullAdder FA_0_5_12_25(S_0_5_12_25, C_0_5_12_25, P_12_13, P_13_12, P_14_11);
	fullAdder FA_0_5_12_26(S_0_5_12_26, C_0_5_12_26, P_12_14, P_13_13, P_14_12);
	fullAdder FA_0_5_12_27(S_0_5_12_27, C_0_5_12_27, P_12_15, P_13_14, P_14_13);
	halfAdder HA_0_5_12_28(S_0_5_12_28, C_0_5_12_28, P_13_15, P_14_14);
 /************************** Height - 1 ********************************/ 
 /************************** Layer - 0 ********************************/ 
	halfAdder HA_1_1_0_2(S_1_1_0_2, C_1_1_0_2, S_0_1_0_2, C_0_1_0_1);
	fullAdder FA_1_1_0_3(S_1_1_0_3, C_1_1_0_3, S_0_1_0_3, C_0_1_0_2, P_3_0);
	fullAdder FA_1_1_0_4(S_1_1_0_4, C_1_1_0_4, S_0_1_0_4, C_0_1_0_3, S_0_2_3_4);
	fullAdder FA_1_1_0_5(S_1_1_0_5, C_1_1_0_5, S_0_1_0_5, C_0_1_0_4, S_0_2_3_5);
	fullAdder FA_1_1_0_6(S_1_1_0_6, C_1_1_0_6, S_0_1_0_6, C_0_1_0_5, S_0_2_3_6);
	fullAdder FA_1_1_0_7(S_1_1_0_7, C_1_1_0_7, S_0_1_0_7, C_0_1_0_6, S_0_2_3_7);
	fullAdder FA_1_1_0_8(S_1_1_0_8, C_1_1_0_8, S_0_1_0_8, C_0_1_0_7, S_0_2_3_8);
	fullAdder FA_1_1_0_9(S_1_1_0_9, C_1_1_0_9, S_0_1_0_9, C_0_1_0_8, S_0_2_3_9);
	fullAdder FA_1_1_0_10(S_1_1_0_10, C_1_1_0_10, S_0_1_0_10, C_0_1_0_9, S_0_2_3_10);
	fullAdder FA_1_1_0_11(S_1_1_0_11, C_1_1_0_11, S_0_1_0_11, C_0_1_0_10, S_0_2_3_11);
	fullAdder FA_1_1_0_12(S_1_1_0_12, C_1_1_0_12, S_0_1_0_12, C_0_1_0_11, S_0_2_3_12);
	fullAdder FA_1_1_0_13(S_1_1_0_13, C_1_1_0_13, S_0_1_0_13, C_0_1_0_12, S_0_2_3_13);
	fullAdder FA_1_1_0_14(S_1_1_0_14, C_1_1_0_14, S_0_1_0_14, C_0_1_0_13, S_0_2_3_14);
	fullAdder FA_1_1_0_15(S_1_1_0_15, C_1_1_0_15, S_0_1_0_15, C_0_1_0_14, S_0_2_3_15);
	fullAdder FA_1_1_0_16(S_1_1_0_16, C_1_1_0_16, S_0_1_0_16, C_0_1_0_15, S_0_2_3_16);
	fullAdder FA_1_1_0_17(S_1_1_0_17, C_1_1_0_17, P_2_15, C_0_1_0_16, S_0_2_3_17);
 /************************** Layer - 3 ********************************/ 
	halfAdder HA_1_2_3_6(S_1_2_3_6, C_1_2_3_6, C_0_2_3_5, P_6_0);
	halfAdder HA_1_2_3_7(S_1_2_3_7, C_1_2_3_7, C_0_2_3_6, S_0_3_6_7);
	fullAdder FA_1_2_3_8(S_1_2_3_8, C_1_2_3_8, C_0_2_3_7, S_0_3_6_8, C_0_3_6_7);
	fullAdder FA_1_2_3_9(S_1_2_3_9, C_1_2_3_9, C_0_2_3_8, S_0_3_6_9, C_0_3_6_8);
	fullAdder FA_1_2_3_10(S_1_2_3_10, C_1_2_3_10, C_0_2_3_9, S_0_3_6_10, C_0_3_6_9);
	fullAdder FA_1_2_3_11(S_1_2_3_11, C_1_2_3_11, C_0_2_3_10, S_0_3_6_11, C_0_3_6_10);
	fullAdder FA_1_2_3_12(S_1_2_3_12, C_1_2_3_12, C_0_2_3_11, S_0_3_6_12, C_0_3_6_11);
	fullAdder FA_1_2_3_13(S_1_2_3_13, C_1_2_3_13, C_0_2_3_12, S_0_3_6_13, C_0_3_6_12);
	fullAdder FA_1_2_3_14(S_1_2_3_14, C_1_2_3_14, C_0_2_3_13, S_0_3_6_14, C_0_3_6_13);
	fullAdder FA_1_2_3_15(S_1_2_3_15, C_1_2_3_15, C_0_2_3_14, S_0_3_6_15, C_0_3_6_14);
	fullAdder FA_1_2_3_16(S_1_2_3_16, C_1_2_3_16, C_0_2_3_15, S_0_3_6_16, C_0_3_6_15);
	fullAdder FA_1_2_3_17(S_1_2_3_17, C_1_2_3_17, C_0_2_3_16, S_0_3_6_17, C_0_3_6_16);
	fullAdder FA_1_2_3_18(S_1_2_3_18, C_1_2_3_18, C_0_2_3_17, S_0_3_6_18, C_0_3_6_17);
	fullAdder FA_1_2_3_19(S_1_2_3_19, C_1_2_3_19, C_0_2_3_18, S_0_3_6_19, C_0_3_6_18);
	fullAdder FA_1_2_3_20(S_1_2_3_20, C_1_2_3_20, C_0_2_3_19, S_0_3_6_20, C_0_3_6_19);
	halfAdder HA_1_2_3_21(S_1_2_3_21, C_1_2_3_21, S_0_3_6_21, C_0_3_6_20);
	halfAdder HA_1_2_3_22(S_1_2_3_22, C_1_2_3_22, S_0_3_6_22, C_0_3_6_21);
	halfAdder HA_1_2_3_23(S_1_2_3_23, C_1_2_3_23, P_8_15, C_0_3_6_22);
 /************************** Layer - 6 ********************************/ 
	halfAdder HA_1_3_6_11(S_1_3_6_11, C_1_3_6_11, S_0_4_9_11, C_0_4_9_10);
	fullAdder FA_1_3_6_12(S_1_3_6_12, C_1_3_6_12, S_0_4_9_12, C_0_4_9_11, P_12_0);
	fullAdder FA_1_3_6_13(S_1_3_6_13, C_1_3_6_13, S_0_4_9_13, C_0_4_9_12, S_0_5_12_13);
	fullAdder FA_1_3_6_14(S_1_3_6_14, C_1_3_6_14, S_0_4_9_14, C_0_4_9_13, S_0_5_12_14);
	fullAdder FA_1_3_6_15(S_1_3_6_15, C_1_3_6_15, S_0_4_9_15, C_0_4_9_14, S_0_5_12_15);
	fullAdder FA_1_3_6_16(S_1_3_6_16, C_1_3_6_16, S_0_4_9_16, C_0_4_9_15, S_0_5_12_16);
	fullAdder FA_1_3_6_17(S_1_3_6_17, C_1_3_6_17, S_0_4_9_17, C_0_4_9_16, S_0_5_12_17);
	fullAdder FA_1_3_6_18(S_1_3_6_18, C_1_3_6_18, S_0_4_9_18, C_0_4_9_17, S_0_5_12_18);
	fullAdder FA_1_3_6_19(S_1_3_6_19, C_1_3_6_19, S_0_4_9_19, C_0_4_9_18, S_0_5_12_19);
	fullAdder FA_1_3_6_20(S_1_3_6_20, C_1_3_6_20, S_0_4_9_20, C_0_4_9_19, S_0_5_12_20);
	fullAdder FA_1_3_6_21(S_1_3_6_21, C_1_3_6_21, S_0_4_9_21, C_0_4_9_20, S_0_5_12_21);
	fullAdder FA_1_3_6_22(S_1_3_6_22, C_1_3_6_22, S_0_4_9_22, C_0_4_9_21, S_0_5_12_22);
	fullAdder FA_1_3_6_23(S_1_3_6_23, C_1_3_6_23, S_0_4_9_23, C_0_4_9_22, S_0_5_12_23);
	fullAdder FA_1_3_6_24(S_1_3_6_24, C_1_3_6_24, S_0_4_9_24, C_0_4_9_23, S_0_5_12_24);
	fullAdder FA_1_3_6_25(S_1_3_6_25, C_1_3_6_25, S_0_4_9_25, C_0_4_9_24, S_0_5_12_25);
	fullAdder FA_1_3_6_26(S_1_3_6_26, C_1_3_6_26, P_11_15, C_0_4_9_25, S_0_5_12_26);
 /************************** Height - 2 ********************************/ 
 /************************** Layer - 0 ********************************/ 
	halfAdder HA_2_1_0_3(S_2_1_0_3, C_2_1_0_3, S_1_1_0_3, C_1_1_0_2);
	halfAdder HA_2_1_0_4(S_2_1_0_4, C_2_1_0_4, S_1_1_0_4, C_1_1_0_3);
	fullAdder FA_2_1_0_5(S_2_1_0_5, C_2_1_0_5, S_1_1_0_5, C_1_1_0_4, C_0_2_3_4);
	fullAdder FA_2_1_0_6(S_2_1_0_6, C_2_1_0_6, S_1_1_0_6, C_1_1_0_5, S_1_2_3_6);
	fullAdder FA_2_1_0_7(S_2_1_0_7, C_2_1_0_7, S_1_1_0_7, C_1_1_0_6, S_1_2_3_7);
	fullAdder FA_2_1_0_8(S_2_1_0_8, C_2_1_0_8, S_1_1_0_8, C_1_1_0_7, S_1_2_3_8);
	fullAdder FA_2_1_0_9(S_2_1_0_9, C_2_1_0_9, S_1_1_0_9, C_1_1_0_8, S_1_2_3_9);
	fullAdder FA_2_1_0_10(S_2_1_0_10, C_2_1_0_10, S_1_1_0_10, C_1_1_0_9, S_1_2_3_10);
	fullAdder FA_2_1_0_11(S_2_1_0_11, C_2_1_0_11, S_1_1_0_11, C_1_1_0_10, S_1_2_3_11);
	fullAdder FA_2_1_0_12(S_2_1_0_12, C_2_1_0_12, S_1_1_0_12, C_1_1_0_11, S_1_2_3_12);
	fullAdder FA_2_1_0_13(S_2_1_0_13, C_2_1_0_13, S_1_1_0_13, C_1_1_0_12, S_1_2_3_13);
	fullAdder FA_2_1_0_14(S_2_1_0_14, C_2_1_0_14, S_1_1_0_14, C_1_1_0_13, S_1_2_3_14);
	fullAdder FA_2_1_0_15(S_2_1_0_15, C_2_1_0_15, S_1_1_0_15, C_1_1_0_14, S_1_2_3_15);
	fullAdder FA_2_1_0_16(S_2_1_0_16, C_2_1_0_16, S_1_1_0_16, C_1_1_0_15, S_1_2_3_16);
	fullAdder FA_2_1_0_17(S_2_1_0_17, C_2_1_0_17, S_1_1_0_17, C_1_1_0_16, S_1_2_3_17);
	fullAdder FA_2_1_0_18(S_2_1_0_18, C_2_1_0_18, S_0_2_3_18, C_1_1_0_17, S_1_2_3_18);
	halfAdder HA_2_1_0_19(S_2_1_0_19, C_2_1_0_19, S_0_2_3_19, S_1_2_3_19);
	halfAdder HA_2_1_0_20(S_2_1_0_20, C_2_1_0_20, P_5_15, S_1_2_3_20);
 /************************** Layer - 3 ********************************/ 
	halfAdder HA_2_2_3_9(S_2_2_3_9, C_2_2_3_9, C_1_2_3_8, P_9_0);
	halfAdder HA_2_2_3_10(S_2_2_3_10, C_2_2_3_10, C_1_2_3_9, S_0_4_9_10);
	halfAdder HA_2_2_3_11(S_2_2_3_11, C_2_2_3_11, C_1_2_3_10, S_1_3_6_11);
	fullAdder FA_2_2_3_12(S_2_2_3_12, C_2_2_3_12, C_1_2_3_11, S_1_3_6_12, C_1_3_6_11);
	fullAdder FA_2_2_3_13(S_2_2_3_13, C_2_2_3_13, C_1_2_3_12, S_1_3_6_13, C_1_3_6_12);
	fullAdder FA_2_2_3_14(S_2_2_3_14, C_2_2_3_14, C_1_2_3_13, S_1_3_6_14, C_1_3_6_13);
	fullAdder FA_2_2_3_15(S_2_2_3_15, C_2_2_3_15, C_1_2_3_14, S_1_3_6_15, C_1_3_6_14);
	fullAdder FA_2_2_3_16(S_2_2_3_16, C_2_2_3_16, C_1_2_3_15, S_1_3_6_16, C_1_3_6_15);
	fullAdder FA_2_2_3_17(S_2_2_3_17, C_2_2_3_17, C_1_2_3_16, S_1_3_6_17, C_1_3_6_16);
	fullAdder FA_2_2_3_18(S_2_2_3_18, C_2_2_3_18, C_1_2_3_17, S_1_3_6_18, C_1_3_6_17);
	fullAdder FA_2_2_3_19(S_2_2_3_19, C_2_2_3_19, C_1_2_3_18, S_1_3_6_19, C_1_3_6_18);
	fullAdder FA_2_2_3_20(S_2_2_3_20, C_2_2_3_20, C_1_2_3_19, S_1_3_6_20, C_1_3_6_19);
	fullAdder FA_2_2_3_21(S_2_2_3_21, C_2_2_3_21, C_1_2_3_20, S_1_3_6_21, C_1_3_6_20);
	fullAdder FA_2_2_3_22(S_2_2_3_22, C_2_2_3_22, C_1_2_3_21, S_1_3_6_22, C_1_3_6_21);
	fullAdder FA_2_2_3_23(S_2_2_3_23, C_2_2_3_23, C_1_2_3_22, S_1_3_6_23, C_1_3_6_22);
	fullAdder FA_2_2_3_24(S_2_2_3_24, C_2_2_3_24, C_1_2_3_23, S_1_3_6_24, C_1_3_6_23);
	halfAdder HA_2_2_3_25(S_2_2_3_25, C_2_2_3_25, S_1_3_6_25, C_1_3_6_24);
	halfAdder HA_2_2_3_26(S_2_2_3_26, C_2_2_3_26, S_1_3_6_26, C_1_3_6_25);
	halfAdder HA_2_2_3_27(S_2_2_3_27, C_2_2_3_27, S_0_5_12_27, C_1_3_6_26);
 /************************** Height - 3 ********************************/ 
 /************************** Layer - 0 ********************************/ 
	halfAdder HA_3_1_0_4(S_3_1_0_4, C_3_1_0_4, S_2_1_0_4, C_2_1_0_3);
	halfAdder HA_3_1_0_5(S_3_1_0_5, C_3_1_0_5, S_2_1_0_5, C_2_1_0_4);
	halfAdder HA_3_1_0_6(S_3_1_0_6, C_3_1_0_6, S_2_1_0_6, C_2_1_0_5);
	fullAdder FA_3_1_0_7(S_3_1_0_7, C_3_1_0_7, S_2_1_0_7, C_2_1_0_6, C_1_2_3_6);
	fullAdder FA_3_1_0_8(S_3_1_0_8, C_3_1_0_8, S_2_1_0_8, C_2_1_0_7, C_1_2_3_7);
	fullAdder FA_3_1_0_9(S_3_1_0_9, C_3_1_0_9, S_2_1_0_9, C_2_1_0_8, S_2_2_3_9);
	fullAdder FA_3_1_0_10(S_3_1_0_10, C_3_1_0_10, S_2_1_0_10, C_2_1_0_9, S_2_2_3_10);
	fullAdder FA_3_1_0_11(S_3_1_0_11, C_3_1_0_11, S_2_1_0_11, C_2_1_0_10, S_2_2_3_11);
	fullAdder FA_3_1_0_12(S_3_1_0_12, C_3_1_0_12, S_2_1_0_12, C_2_1_0_11, S_2_2_3_12);
	fullAdder FA_3_1_0_13(S_3_1_0_13, C_3_1_0_13, S_2_1_0_13, C_2_1_0_12, S_2_2_3_13);
	fullAdder FA_3_1_0_14(S_3_1_0_14, C_3_1_0_14, S_2_1_0_14, C_2_1_0_13, S_2_2_3_14);
	fullAdder FA_3_1_0_15(S_3_1_0_15, C_3_1_0_15, S_2_1_0_15, C_2_1_0_14, S_2_2_3_15);
	fullAdder FA_3_1_0_16(S_3_1_0_16, C_3_1_0_16, S_2_1_0_16, C_2_1_0_15, S_2_2_3_16);
	fullAdder FA_3_1_0_17(S_3_1_0_17, C_3_1_0_17, S_2_1_0_17, C_2_1_0_16, S_2_2_3_17);
	fullAdder FA_3_1_0_18(S_3_1_0_18, C_3_1_0_18, S_2_1_0_18, C_2_1_0_17, S_2_2_3_18);
	fullAdder FA_3_1_0_19(S_3_1_0_19, C_3_1_0_19, S_2_1_0_19, C_2_1_0_18, S_2_2_3_19);
	fullAdder FA_3_1_0_20(S_3_1_0_20, C_3_1_0_20, S_2_1_0_20, C_2_1_0_19, S_2_2_3_20);
	fullAdder FA_3_1_0_21(S_3_1_0_21, C_3_1_0_21, S_1_2_3_21, C_2_1_0_20, S_2_2_3_21);
	halfAdder HA_3_1_0_22(S_3_1_0_22, C_3_1_0_22, S_1_2_3_22, S_2_2_3_22);
	halfAdder HA_3_1_0_23(S_3_1_0_23, C_3_1_0_23, S_1_2_3_23, S_2_2_3_23);
 /************************** Layer - 3 ********************************/ 
	halfAdder HA_3_2_3_14(S_3_2_3_14, C_3_2_3_14, C_2_2_3_13, C_0_5_12_13);
	fullAdder FA_3_2_3_15(S_3_2_3_15, C_3_2_3_15, C_2_2_3_14, C_0_5_12_14, P_15_0);
	fullAdder FA_3_2_3_16(S_3_2_3_16, C_3_2_3_16, C_2_2_3_15, C_0_5_12_15, P_15_1);
	fullAdder FA_3_2_3_17(S_3_2_3_17, C_3_2_3_17, C_2_2_3_16, C_0_5_12_16, P_15_2);
	fullAdder FA_3_2_3_18(S_3_2_3_18, C_3_2_3_18, C_2_2_3_17, C_0_5_12_17, P_15_3);
	fullAdder FA_3_2_3_19(S_3_2_3_19, C_3_2_3_19, C_2_2_3_18, C_0_5_12_18, P_15_4);
	fullAdder FA_3_2_3_20(S_3_2_3_20, C_3_2_3_20, C_2_2_3_19, C_0_5_12_19, P_15_5);
	fullAdder FA_3_2_3_21(S_3_2_3_21, C_3_2_3_21, C_2_2_3_20, C_0_5_12_20, P_15_6);
	fullAdder FA_3_2_3_22(S_3_2_3_22, C_3_2_3_22, C_2_2_3_21, C_0_5_12_21, P_15_7);
	fullAdder FA_3_2_3_23(S_3_2_3_23, C_3_2_3_23, C_2_2_3_22, C_0_5_12_22, P_15_8);
	fullAdder FA_3_2_3_24(S_3_2_3_24, C_3_2_3_24, C_2_2_3_23, C_0_5_12_23, P_15_9);
	fullAdder FA_3_2_3_25(S_3_2_3_25, C_3_2_3_25, C_2_2_3_24, C_0_5_12_24, P_15_10);
	fullAdder FA_3_2_3_26(S_3_2_3_26, C_3_2_3_26, C_2_2_3_25, C_0_5_12_25, P_15_11);
	fullAdder FA_3_2_3_27(S_3_2_3_27, C_3_2_3_27, C_2_2_3_26, C_0_5_12_26, P_15_12);
	fullAdder FA_3_2_3_28(S_3_2_3_28, C_3_2_3_28, C_2_2_3_27, C_0_5_12_27, P_15_13);
	halfAdder HA_3_2_3_29(S_3_2_3_29, C_3_2_3_29, C_0_5_12_28, P_15_14);
 /************************** Height - 4 ********************************/ 
 /************************** Layer - 0 ********************************/ 
	halfAdder HA_4_1_0_5(S_4_1_0_5, C_4_1_0_5, S_3_1_0_5, C_3_1_0_4);
	halfAdder HA_4_1_0_6(S_4_1_0_6, C_4_1_0_6, S_3_1_0_6, C_3_1_0_5);
	halfAdder HA_4_1_0_7(S_4_1_0_7, C_4_1_0_7, S_3_1_0_7, C_3_1_0_6);
	halfAdder HA_4_1_0_8(S_4_1_0_8, C_4_1_0_8, S_3_1_0_8, C_3_1_0_7);
	halfAdder HA_4_1_0_9(S_4_1_0_9, C_4_1_0_9, S_3_1_0_9, C_3_1_0_8);
	fullAdder FA_4_1_0_10(S_4_1_0_10, C_4_1_0_10, S_3_1_0_10, C_3_1_0_9, C_2_2_3_9);
	fullAdder FA_4_1_0_11(S_4_1_0_11, C_4_1_0_11, S_3_1_0_11, C_3_1_0_10, C_2_2_3_10);
	fullAdder FA_4_1_0_12(S_4_1_0_12, C_4_1_0_12, S_3_1_0_12, C_3_1_0_11, C_2_2_3_11);
	fullAdder FA_4_1_0_13(S_4_1_0_13, C_4_1_0_13, S_3_1_0_13, C_3_1_0_12, C_2_2_3_12);
	fullAdder FA_4_1_0_14(S_4_1_0_14, C_4_1_0_14, S_3_1_0_14, C_3_1_0_13, S_3_2_3_14);
	fullAdder FA_4_1_0_15(S_4_1_0_15, C_4_1_0_15, S_3_1_0_15, C_3_1_0_14, S_3_2_3_15);
	fullAdder FA_4_1_0_16(S_4_1_0_16, C_4_1_0_16, S_3_1_0_16, C_3_1_0_15, S_3_2_3_16);
	fullAdder FA_4_1_0_17(S_4_1_0_17, C_4_1_0_17, S_3_1_0_17, C_3_1_0_16, S_3_2_3_17);
	fullAdder FA_4_1_0_18(S_4_1_0_18, C_4_1_0_18, S_3_1_0_18, C_3_1_0_17, S_3_2_3_18);
	fullAdder FA_4_1_0_19(S_4_1_0_19, C_4_1_0_19, S_3_1_0_19, C_3_1_0_18, S_3_2_3_19);
	fullAdder FA_4_1_0_20(S_4_1_0_20, C_4_1_0_20, S_3_1_0_20, C_3_1_0_19, S_3_2_3_20);
	fullAdder FA_4_1_0_21(S_4_1_0_21, C_4_1_0_21, S_3_1_0_21, C_3_1_0_20, S_3_2_3_21);
	fullAdder FA_4_1_0_22(S_4_1_0_22, C_4_1_0_22, S_3_1_0_22, C_3_1_0_21, S_3_2_3_22);
	fullAdder FA_4_1_0_23(S_4_1_0_23, C_4_1_0_23, S_3_1_0_23, C_3_1_0_22, S_3_2_3_23);
	fullAdder FA_4_1_0_24(S_4_1_0_24, C_4_1_0_24, S_2_2_3_24, C_3_1_0_23, S_3_2_3_24);
	halfAdder HA_4_1_0_25(S_4_1_0_25, C_4_1_0_25, S_2_2_3_25, S_3_2_3_25);
	halfAdder HA_4_1_0_26(S_4_1_0_26, C_4_1_0_26, S_2_2_3_26, S_3_2_3_26);
	halfAdder HA_4_1_0_27(S_4_1_0_27, C_4_1_0_27, S_2_2_3_27, S_3_2_3_27);
	halfAdder HA_4_1_0_28(S_4_1_0_28, C_4_1_0_28, S_0_5_12_28, S_3_2_3_28);
	halfAdder HA_4_1_0_29(S_4_1_0_29, C_4_1_0_29, P_14_15, S_3_2_3_29);
 /************************** Height - 5 ********************************/ 
 /************************** Layer - 0 ********************************/ 
	halfAdder HA_5_1_0_6(S_5_1_0_6, C_5_1_0_6, S_4_1_0_6, C_4_1_0_5);
	halfAdder HA_5_1_0_7(S_5_1_0_7, C_5_1_0_7, S_4_1_0_7, C_4_1_0_6);
	halfAdder HA_5_1_0_8(S_5_1_0_8, C_5_1_0_8, S_4_1_0_8, C_4_1_0_7);
	halfAdder HA_5_1_0_9(S_5_1_0_9, C_5_1_0_9, S_4_1_0_9, C_4_1_0_8);
	halfAdder HA_5_1_0_10(S_5_1_0_10, C_5_1_0_10, S_4_1_0_10, C_4_1_0_9);
	halfAdder HA_5_1_0_11(S_5_1_0_11, C_5_1_0_11, S_4_1_0_11, C_4_1_0_10);
	halfAdder HA_5_1_0_12(S_5_1_0_12, C_5_1_0_12, S_4_1_0_12, C_4_1_0_11);
	halfAdder HA_5_1_0_13(S_5_1_0_13, C_5_1_0_13, S_4_1_0_13, C_4_1_0_12);
	halfAdder HA_5_1_0_14(S_5_1_0_14, C_5_1_0_14, S_4_1_0_14, C_4_1_0_13);
	fullAdder FA_5_1_0_15(S_5_1_0_15, C_5_1_0_15, S_4_1_0_15, C_4_1_0_14, C_3_2_3_14);
	fullAdder FA_5_1_0_16(S_5_1_0_16, C_5_1_0_16, S_4_1_0_16, C_4_1_0_15, C_3_2_3_15);
	fullAdder FA_5_1_0_17(S_5_1_0_17, C_5_1_0_17, S_4_1_0_17, C_4_1_0_16, C_3_2_3_16);
	fullAdder FA_5_1_0_18(S_5_1_0_18, C_5_1_0_18, S_4_1_0_18, C_4_1_0_17, C_3_2_3_17);
	fullAdder FA_5_1_0_19(S_5_1_0_19, C_5_1_0_19, S_4_1_0_19, C_4_1_0_18, C_3_2_3_18);
	fullAdder FA_5_1_0_20(S_5_1_0_20, C_5_1_0_20, S_4_1_0_20, C_4_1_0_19, C_3_2_3_19);
	fullAdder FA_5_1_0_21(S_5_1_0_21, C_5_1_0_21, S_4_1_0_21, C_4_1_0_20, C_3_2_3_20);
	fullAdder FA_5_1_0_22(S_5_1_0_22, C_5_1_0_22, S_4_1_0_22, C_4_1_0_21, C_3_2_3_21);
	fullAdder FA_5_1_0_23(S_5_1_0_23, C_5_1_0_23, S_4_1_0_23, C_4_1_0_22, C_3_2_3_22);
	fullAdder FA_5_1_0_24(S_5_1_0_24, C_5_1_0_24, S_4_1_0_24, C_4_1_0_23, C_3_2_3_23);
	fullAdder FA_5_1_0_25(S_5_1_0_25, C_5_1_0_25, S_4_1_0_25, C_4_1_0_24, C_3_2_3_24);
	fullAdder FA_5_1_0_26(S_5_1_0_26, C_5_1_0_26, S_4_1_0_26, C_4_1_0_25, C_3_2_3_25);
	fullAdder FA_5_1_0_27(S_5_1_0_27, C_5_1_0_27, S_4_1_0_27, C_4_1_0_26, C_3_2_3_26);
	fullAdder FA_5_1_0_28(S_5_1_0_28, C_5_1_0_28, S_4_1_0_28, C_4_1_0_27, C_3_2_3_27);
	fullAdder FA_5_1_0_29(S_5_1_0_29, C_5_1_0_29, S_4_1_0_29, C_4_1_0_28, C_3_2_3_28);
	fullAdder FA_5_1_0_30(S_5_1_0_30, C_5_1_0_30, P_15_15, C_4_1_0_29, C_3_2_3_29);


	wire [24:0] in1 = {1'b0, S_5_1_0_30, S_5_1_0_29, S_5_1_0_28, S_5_1_0_27, S_5_1_0_26, S_5_1_0_25, S_5_1_0_24, S_5_1_0_23, S_5_1_0_22, S_5_1_0_21, S_5_1_0_20, S_5_1_0_19, S_5_1_0_18, S_5_1_0_17, S_5_1_0_16, S_5_1_0_15, S_5_1_0_14, S_5_1_0_13, S_5_1_0_12, S_5_1_0_11, S_5_1_0_10, S_5_1_0_9, S_5_1_0_8, S_5_1_0_7};
	wire [24:0] in2 = {C_5_1_0_30, C_5_1_0_29, C_5_1_0_28, C_5_1_0_27, C_5_1_0_26, C_5_1_0_25, C_5_1_0_24, C_5_1_0_23, C_5_1_0_22, C_5_1_0_21, C_5_1_0_20, C_5_1_0_19, C_5_1_0_18, C_5_1_0_17, C_5_1_0_16, C_5_1_0_15, C_5_1_0_14, C_5_1_0_13, C_5_1_0_12, C_5_1_0_11, C_5_1_0_10, C_5_1_0_9, C_5_1_0_8, C_5_1_0_7, C_5_1_0_6};
	wire [24:0] sum;
	assign sum = in1 + in2;
	assign out = {sum, S_5_1_0_6, S_4_1_0_5, S_3_1_0_4, S_2_1_0_3, S_1_1_0_2, S_0_1_0_1, P_0_0};

	endmodule
	